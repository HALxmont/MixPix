magic
tech sky130A
magscale 1 2
timestamp 1668518072
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 410518 700408 410524 700460
rect 410576 700448 410582 700460
rect 429838 700448 429844 700460
rect 410576 700420 429844 700448
rect 410576 700408 410582 700420
rect 429838 700408 429844 700420
rect 429896 700408 429902 700460
rect 409138 700340 409144 700392
rect 409196 700380 409202 700392
rect 494790 700380 494796 700392
rect 409196 700352 494796 700380
rect 409196 700340 409202 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 364978 700272 364984 700324
rect 365036 700312 365042 700324
rect 374638 700312 374644 700324
rect 365036 700284 374644 700312
rect 365036 700272 365042 700284
rect 374638 700272 374644 700284
rect 374696 700272 374702 700324
rect 407758 700272 407764 700324
rect 407816 700312 407822 700324
rect 559650 700312 559656 700324
rect 407816 700284 559656 700312
rect 407816 700272 407822 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 332502 699796 332508 699848
rect 332560 699836 332566 699848
rect 334618 699836 334624 699848
rect 332560 699808 334624 699836
rect 332560 699796 332566 699808
rect 334618 699796 334624 699808
rect 334676 699796 334682 699848
rect 150434 699660 150440 699712
rect 150492 699700 150498 699712
rect 154114 699700 154120 699712
rect 150492 699672 154120 699700
rect 150492 699660 150498 699672
rect 154114 699660 154120 699672
rect 154172 699660 154178 699712
rect 195974 699660 195980 699712
rect 196032 699700 196038 699712
rect 202782 699700 202788 699712
rect 196032 699672 202788 699700
rect 196032 699660 196038 699672
rect 202782 699660 202788 699672
rect 202840 699660 202846 699712
rect 231854 699660 231860 699712
rect 231912 699700 231918 699712
rect 235166 699700 235172 699712
rect 231912 699672 235172 699700
rect 231912 699660 231918 699672
rect 235166 699660 235172 699672
rect 235224 699660 235230 699712
rect 348786 699660 348792 699712
rect 348844 699700 348850 699712
rect 350534 699700 350540 699712
rect 348844 699672 350540 699700
rect 348844 699660 348850 699672
rect 350534 699660 350540 699672
rect 350592 699660 350598 699712
rect 281534 698300 281540 698352
rect 281592 698340 281598 698352
rect 283834 698340 283840 698352
rect 281592 698312 283840 698340
rect 281592 698300 281598 698312
rect 283834 698300 283840 698312
rect 283892 698300 283898 698352
rect 300118 698096 300124 698148
rect 300176 698136 300182 698148
rect 302878 698136 302884 698148
rect 300176 698108 302884 698136
rect 300176 698096 300182 698108
rect 302878 698096 302884 698108
rect 302936 698096 302942 698148
rect 350534 698028 350540 698080
rect 350592 698068 350598 698080
rect 353938 698068 353944 698080
rect 350592 698040 353944 698068
rect 350592 698028 350598 698040
rect 353938 698028 353944 698040
rect 353996 698028 354002 698080
rect 229738 695240 229744 695292
rect 229796 695280 229802 695292
rect 231854 695280 231860 695292
rect 229796 695252 231860 695280
rect 229796 695240 229802 695252
rect 231854 695240 231860 695252
rect 231912 695240 231918 695292
rect 280798 694968 280804 695020
rect 280856 695008 280862 695020
rect 281534 695008 281540 695020
rect 280856 694980 281540 695008
rect 280856 694968 280862 694980
rect 281534 694968 281540 694980
rect 281592 694968 281598 695020
rect 189074 694764 189080 694816
rect 189132 694804 189138 694816
rect 195974 694804 195980 694816
rect 189132 694776 195980 694804
rect 189132 694764 189138 694776
rect 195974 694764 195980 694776
rect 196032 694764 196038 694816
rect 258074 694220 258080 694272
rect 258132 694260 258138 694272
rect 267642 694260 267648 694272
rect 258132 694232 267648 694260
rect 258132 694220 258138 694232
rect 267642 694220 267648 694232
rect 267700 694220 267706 694272
rect 149790 693472 149796 693524
rect 149848 693512 149854 693524
rect 150434 693512 150440 693524
rect 149848 693484 150440 693512
rect 149848 693472 149854 693484
rect 150434 693472 150440 693484
rect 150492 693472 150498 693524
rect 302878 692044 302884 692096
rect 302936 692084 302942 692096
rect 313918 692084 313924 692096
rect 302936 692056 313924 692084
rect 302936 692044 302942 692056
rect 313918 692044 313924 692056
rect 313976 692044 313982 692096
rect 374638 691092 374644 691144
rect 374696 691132 374702 691144
rect 377398 691132 377404 691144
rect 374696 691104 377404 691132
rect 374696 691092 374702 691104
rect 377398 691092 377404 691104
rect 377456 691092 377462 691144
rect 247678 689256 247684 689308
rect 247736 689296 247742 689308
rect 258074 689296 258080 689308
rect 247736 689268 258080 689296
rect 247736 689256 247742 689268
rect 258074 689256 258080 689268
rect 258132 689256 258138 689308
rect 181438 688644 181444 688696
rect 181496 688684 181502 688696
rect 189074 688684 189080 688696
rect 181496 688656 189080 688684
rect 181496 688644 181502 688656
rect 189074 688644 189080 688656
rect 189132 688644 189138 688696
rect 206278 687896 206284 687948
rect 206336 687936 206342 687948
rect 218054 687936 218060 687948
rect 206336 687908 218060 687936
rect 206336 687896 206342 687908
rect 218054 687896 218060 687908
rect 218112 687896 218118 687948
rect 148318 687488 148324 687540
rect 148376 687528 148382 687540
rect 149790 687528 149796 687540
rect 148376 687500 149796 687528
rect 148376 687488 148382 687500
rect 149790 687488 149796 687500
rect 149848 687488 149854 687540
rect 334618 686468 334624 686520
rect 334676 686508 334682 686520
rect 349798 686508 349804 686520
rect 334676 686480 349804 686508
rect 334676 686468 334682 686480
rect 349798 686468 349804 686480
rect 349856 686468 349862 686520
rect 221458 685108 221464 685160
rect 221516 685148 221522 685160
rect 229738 685148 229744 685160
rect 221516 685120 229744 685148
rect 221516 685108 221522 685120
rect 229738 685108 229744 685120
rect 229796 685108 229802 685160
rect 353938 683748 353944 683800
rect 353996 683788 354002 683800
rect 358354 683788 358360 683800
rect 353996 683760 358360 683788
rect 353996 683748 354002 683760
rect 358354 683748 358360 683760
rect 358412 683748 358418 683800
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 313918 682388 313924 682440
rect 313976 682428 313982 682440
rect 333238 682428 333244 682440
rect 313976 682400 333244 682428
rect 313976 682388 313982 682400
rect 333238 682388 333244 682400
rect 333296 682388 333302 682440
rect 204254 681708 204260 681760
rect 204312 681748 204318 681760
rect 206278 681748 206284 681760
rect 204312 681720 206284 681748
rect 204312 681708 204318 681720
rect 206278 681708 206284 681720
rect 206336 681708 206342 681760
rect 148318 679028 148324 679040
rect 146312 679000 148324 679028
rect 144178 678920 144184 678972
rect 144236 678960 144242 678972
rect 146312 678960 146340 679000
rect 148318 678988 148324 679000
rect 148376 678988 148382 679040
rect 144236 678932 146340 678960
rect 144236 678920 144242 678932
rect 358354 678444 358360 678496
rect 358412 678484 358418 678496
rect 360838 678484 360844 678496
rect 358412 678456 360844 678484
rect 358412 678444 358418 678456
rect 360838 678444 360844 678456
rect 360896 678444 360902 678496
rect 377398 678240 377404 678292
rect 377456 678280 377462 678292
rect 396442 678280 396448 678292
rect 377456 678252 396448 678280
rect 377456 678240 377462 678252
rect 396442 678240 396448 678252
rect 396500 678240 396506 678292
rect 202138 677016 202144 677068
rect 202196 677056 202202 677068
rect 204254 677056 204260 677068
rect 202196 677028 204260 677056
rect 202196 677016 202202 677028
rect 204254 677016 204260 677028
rect 204312 677016 204318 677068
rect 166994 671304 167000 671356
rect 167052 671344 167058 671356
rect 181438 671344 181444 671356
rect 167052 671316 181444 671344
rect 167052 671304 167058 671316
rect 181438 671304 181444 671316
rect 181496 671304 181502 671356
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 406378 670692 406384 670744
rect 406436 670732 406442 670744
rect 580166 670732 580172 670744
rect 406436 670704 580172 670732
rect 406436 670692 406442 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 215938 668584 215944 668636
rect 215996 668624 216002 668636
rect 221458 668624 221464 668636
rect 215996 668596 221464 668624
rect 215996 668584 216002 668596
rect 221458 668584 221464 668596
rect 221516 668584 221522 668636
rect 360838 668584 360844 668636
rect 360896 668624 360902 668636
rect 363598 668624 363604 668636
rect 360896 668596 363604 668624
rect 360896 668584 360902 668596
rect 363598 668584 363604 668596
rect 363656 668584 363662 668636
rect 160738 667156 160744 667208
rect 160796 667196 160802 667208
rect 166994 667196 167000 667208
rect 160796 667168 167000 667196
rect 160796 667156 160802 667168
rect 166994 667156 167000 667168
rect 167052 667156 167058 667208
rect 200114 666340 200120 666392
rect 200172 666380 200178 666392
rect 202138 666380 202144 666392
rect 200172 666352 202144 666380
rect 200172 666340 200178 666352
rect 202138 666340 202144 666352
rect 202196 666340 202202 666392
rect 279418 665116 279424 665168
rect 279476 665156 279482 665168
rect 280798 665156 280804 665168
rect 279476 665128 280804 665156
rect 279476 665116 279482 665128
rect 280798 665116 280804 665128
rect 280856 665116 280862 665168
rect 363598 663008 363604 663060
rect 363656 663048 363662 663060
rect 369118 663048 369124 663060
rect 363656 663020 369124 663048
rect 363656 663008 363662 663020
rect 369118 663008 369124 663020
rect 369176 663008 369182 663060
rect 141418 662396 141424 662448
rect 141476 662436 141482 662448
rect 144178 662436 144184 662448
rect 141476 662408 144184 662436
rect 141476 662396 141482 662408
rect 144178 662396 144184 662408
rect 144236 662396 144242 662448
rect 153838 661036 153844 661088
rect 153896 661076 153902 661088
rect 160738 661076 160744 661088
rect 153896 661048 160744 661076
rect 153896 661036 153902 661048
rect 160738 661036 160744 661048
rect 160796 661036 160802 661088
rect 369118 660288 369124 660340
rect 369176 660328 369182 660340
rect 387334 660328 387340 660340
rect 369176 660300 387340 660328
rect 369176 660288 369182 660300
rect 387334 660288 387340 660300
rect 387392 660288 387398 660340
rect 195146 659200 195152 659252
rect 195204 659240 195210 659252
rect 200114 659240 200120 659252
rect 195204 659212 200120 659240
rect 195204 659200 195210 659212
rect 200114 659200 200120 659212
rect 200172 659200 200178 659252
rect 241974 658928 241980 658980
rect 242032 658968 242038 658980
rect 247678 658968 247684 658980
rect 242032 658940 247684 658968
rect 242032 658928 242038 658940
rect 247678 658928 247684 658940
rect 247736 658928 247742 658980
rect 349798 658180 349804 658232
rect 349856 658220 349862 658232
rect 355778 658220 355784 658232
rect 349856 658192 355784 658220
rect 349856 658180 349862 658192
rect 355778 658180 355784 658192
rect 355836 658180 355842 658232
rect 387334 658180 387340 658232
rect 387392 658220 387398 658232
rect 393958 658220 393964 658232
rect 387392 658192 393964 658220
rect 387392 658180 387398 658192
rect 393958 658180 393964 658192
rect 394016 658180 394022 658232
rect 235258 656140 235264 656192
rect 235316 656180 235322 656192
rect 241974 656180 241980 656192
rect 235316 656152 241980 656180
rect 235316 656140 235322 656152
rect 241974 656140 241980 656152
rect 242032 656140 242038 656192
rect 274634 655528 274640 655580
rect 274692 655568 274698 655580
rect 279418 655568 279424 655580
rect 274692 655540 279424 655568
rect 274692 655528 274698 655540
rect 279418 655528 279424 655540
rect 279476 655528 279482 655580
rect 355778 655460 355784 655512
rect 355836 655500 355842 655512
rect 358722 655500 358728 655512
rect 355836 655472 358728 655500
rect 355836 655460 355842 655472
rect 358722 655460 358728 655472
rect 358780 655460 358786 655512
rect 185578 654780 185584 654832
rect 185636 654820 185642 654832
rect 195146 654820 195152 654832
rect 185636 654792 195152 654820
rect 185636 654780 185642 654792
rect 195146 654780 195152 654792
rect 195204 654780 195210 654832
rect 273898 652740 273904 652792
rect 273956 652780 273962 652792
rect 274634 652780 274640 652792
rect 273956 652752 274640 652780
rect 273956 652740 273962 652752
rect 274634 652740 274640 652752
rect 274692 652740 274698 652792
rect 146938 651992 146944 652044
rect 146996 652032 147002 652044
rect 153838 652032 153844 652044
rect 146996 652004 153844 652032
rect 146996 651992 147002 652004
rect 153838 651992 153844 652004
rect 153896 651992 153902 652044
rect 358722 650632 358728 650684
rect 358780 650672 358786 650684
rect 369118 650672 369124 650684
rect 358780 650644 369124 650672
rect 358780 650632 358786 650644
rect 369118 650632 369124 650644
rect 369176 650632 369182 650684
rect 393958 649884 393964 649936
rect 394016 649924 394022 649936
rect 395338 649924 395344 649936
rect 394016 649896 395344 649924
rect 394016 649884 394022 649896
rect 395338 649884 395344 649896
rect 395396 649884 395402 649936
rect 203518 647844 203524 647896
rect 203576 647884 203582 647896
rect 215938 647884 215944 647896
rect 203576 647856 215944 647884
rect 203576 647844 203582 647856
rect 215938 647844 215944 647856
rect 215996 647844 216002 647896
rect 395338 647164 395344 647216
rect 395396 647204 395402 647216
rect 396534 647204 396540 647216
rect 395396 647176 396540 647204
rect 395396 647164 395402 647176
rect 396534 647164 396540 647176
rect 396592 647164 396598 647216
rect 333238 643696 333244 643748
rect 333296 643736 333302 643748
rect 353938 643736 353944 643748
rect 333296 643708 353944 643736
rect 333296 643696 333302 643708
rect 353938 643696 353944 643708
rect 353996 643696 354002 643748
rect 396718 643084 396724 643136
rect 396776 643124 396782 643136
rect 580166 643124 580172 643136
rect 396776 643096 580172 643124
rect 396776 643084 396782 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 144178 641724 144184 641776
rect 144236 641764 144242 641776
rect 146938 641764 146944 641776
rect 144236 641736 146944 641764
rect 144236 641724 144242 641736
rect 146938 641724 146944 641736
rect 146996 641724 147002 641776
rect 369118 640500 369124 640552
rect 369176 640540 369182 640552
rect 371878 640540 371884 640552
rect 369176 640512 371884 640540
rect 369176 640500 369182 640512
rect 371878 640500 371884 640512
rect 371936 640500 371942 640552
rect 232498 639412 232504 639464
rect 232556 639452 232562 639464
rect 235258 639452 235264 639464
rect 232556 639424 235264 639452
rect 232556 639412 232562 639424
rect 235258 639412 235264 639424
rect 235316 639412 235322 639464
rect 140038 638188 140044 638240
rect 140096 638228 140102 638240
rect 141418 638228 141424 638240
rect 140096 638200 141424 638228
rect 140096 638188 140102 638200
rect 141418 638188 141424 638200
rect 141476 638188 141482 638240
rect 196618 635468 196624 635520
rect 196676 635508 196682 635520
rect 203518 635508 203524 635520
rect 196676 635480 203524 635508
rect 196676 635468 196682 635480
rect 203518 635468 203524 635480
rect 203576 635468 203582 635520
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4890 632108 4896 632120
rect 2832 632080 4896 632108
rect 2832 632068 2838 632080
rect 4890 632068 4896 632080
rect 4948 632068 4954 632120
rect 184198 632068 184204 632120
rect 184256 632108 184262 632120
rect 185578 632108 185584 632120
rect 184256 632080 185584 632108
rect 184256 632068 184262 632080
rect 185578 632068 185584 632080
rect 185636 632068 185642 632120
rect 272610 632068 272616 632120
rect 272668 632108 272674 632120
rect 273898 632108 273904 632120
rect 272668 632080 273904 632108
rect 272668 632068 272674 632080
rect 273898 632068 273904 632080
rect 273956 632068 273962 632120
rect 271138 629688 271144 629740
rect 271196 629728 271202 629740
rect 272610 629728 272616 629740
rect 271196 629700 272616 629728
rect 271196 629688 271202 629700
rect 272610 629688 272616 629700
rect 272668 629688 272674 629740
rect 140038 627960 140044 627972
rect 138032 627932 140044 627960
rect 136358 627852 136364 627904
rect 136416 627892 136422 627904
rect 138032 627892 138060 627932
rect 140038 627920 140044 627932
rect 140096 627920 140102 627972
rect 136416 627864 138060 627892
rect 136416 627852 136422 627864
rect 353938 625812 353944 625864
rect 353996 625852 354002 625864
rect 395338 625852 395344 625864
rect 353996 625824 395344 625852
rect 353996 625812 354002 625824
rect 395338 625812 395344 625824
rect 395396 625812 395402 625864
rect 134518 620304 134524 620356
rect 134576 620344 134582 620356
rect 136358 620344 136364 620356
rect 134576 620316 136364 620344
rect 134576 620304 134582 620316
rect 136358 620304 136364 620316
rect 136416 620304 136422 620356
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 19978 618304 19984 618316
rect 3568 618276 19984 618304
rect 3568 618264 3574 618276
rect 19978 618264 19984 618276
rect 20036 618264 20042 618316
rect 404998 616836 405004 616888
rect 405056 616876 405062 616888
rect 580166 616876 580172 616888
rect 405056 616848 580172 616876
rect 405056 616836 405062 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 269390 616768 269396 616820
rect 269448 616808 269454 616820
rect 271138 616808 271144 616820
rect 269448 616780 271144 616808
rect 269448 616768 269454 616780
rect 271138 616768 271144 616780
rect 271196 616768 271202 616820
rect 126238 608744 126244 608796
rect 126296 608784 126302 608796
rect 134518 608784 134524 608796
rect 126296 608756 134524 608784
rect 126296 608744 126302 608756
rect 134518 608744 134524 608756
rect 134576 608744 134582 608796
rect 268378 608744 268384 608796
rect 268436 608784 268442 608796
rect 269390 608784 269396 608796
rect 268436 608756 269396 608784
rect 268436 608744 268442 608756
rect 269390 608744 269396 608756
rect 269448 608744 269454 608796
rect 182818 603100 182824 603152
rect 182876 603140 182882 603152
rect 184198 603140 184204 603152
rect 182876 603112 184204 603140
rect 182876 603100 182882 603112
rect 184198 603100 184204 603112
rect 184256 603100 184262 603152
rect 137738 597524 137744 597576
rect 137796 597564 137802 597576
rect 144178 597564 144184 597576
rect 137796 597536 144184 597564
rect 137796 597524 137802 597536
rect 144178 597524 144184 597536
rect 144236 597524 144242 597576
rect 264238 593512 264244 593564
rect 264296 593552 264302 593564
rect 268378 593552 268384 593564
rect 264296 593524 268384 593552
rect 264296 593512 264302 593524
rect 268378 593512 268384 593524
rect 268436 593512 268442 593564
rect 133138 592016 133144 592068
rect 133196 592056 133202 592068
rect 137738 592056 137744 592068
rect 133196 592028 137744 592056
rect 133196 592016 133202 592028
rect 137738 592016 137744 592028
rect 137796 592016 137802 592068
rect 120718 591268 120724 591320
rect 120776 591308 120782 591320
rect 126238 591308 126244 591320
rect 120776 591280 126244 591308
rect 120776 591268 120782 591280
rect 126238 591268 126244 591280
rect 126296 591268 126302 591320
rect 371878 591268 371884 591320
rect 371936 591308 371942 591320
rect 384298 591308 384304 591320
rect 371936 591280 384304 591308
rect 371936 591268 371942 591280
rect 384298 591268 384304 591280
rect 384356 591268 384362 591320
rect 229738 590316 229744 590368
rect 229796 590356 229802 590368
rect 232498 590356 232504 590368
rect 229796 590328 232504 590356
rect 229796 590316 229802 590328
rect 232498 590316 232504 590328
rect 232556 590316 232562 590368
rect 119338 585148 119344 585200
rect 119396 585188 119402 585200
rect 120718 585188 120724 585200
rect 119396 585160 120724 585188
rect 119396 585148 119402 585160
rect 120718 585148 120724 585160
rect 120776 585148 120782 585200
rect 262858 585148 262864 585200
rect 262916 585188 262922 585200
rect 264238 585188 264244 585200
rect 262916 585160 264244 585188
rect 262916 585148 262922 585160
rect 264238 585148 264244 585160
rect 264296 585148 264302 585200
rect 384298 583516 384304 583568
rect 384356 583556 384362 583568
rect 390554 583556 390560 583568
rect 384356 583528 390560 583556
rect 384356 583516 384362 583528
rect 390554 583516 390560 583528
rect 390612 583516 390618 583568
rect 207658 581612 207664 581664
rect 207716 581652 207722 581664
rect 229738 581652 229744 581664
rect 207716 581624 229744 581652
rect 207716 581612 207722 581624
rect 229738 581612 229744 581624
rect 229796 581612 229802 581664
rect 3510 579640 3516 579692
rect 3568 579680 3574 579692
rect 10318 579680 10324 579692
rect 3568 579652 10324 579680
rect 3568 579640 3574 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 129734 578212 129740 578264
rect 129792 578252 129798 578264
rect 133138 578252 133144 578264
rect 129792 578224 133144 578252
rect 129792 578212 129798 578224
rect 133138 578212 133144 578224
rect 133196 578212 133202 578264
rect 181438 578144 181444 578196
rect 181496 578184 181502 578196
rect 182818 578184 182824 578196
rect 181496 578156 182824 578184
rect 181496 578144 181502 578156
rect 182818 578144 182824 578156
rect 182876 578144 182882 578196
rect 390554 576852 390560 576904
rect 390612 576892 390618 576904
rect 393958 576892 393964 576904
rect 390612 576864 393964 576892
rect 390612 576852 390618 576864
rect 393958 576852 393964 576864
rect 394016 576852 394022 576904
rect 120718 570596 120724 570648
rect 120776 570636 120782 570648
rect 129734 570636 129740 570648
rect 120776 570608 129740 570636
rect 120776 570596 120782 570608
rect 129734 570596 129740 570608
rect 129792 570596 129798 570648
rect 261478 570596 261484 570648
rect 261536 570636 261542 570648
rect 262858 570636 262864 570648
rect 261536 570608 262864 570636
rect 261536 570596 261542 570608
rect 262858 570596 262864 570608
rect 262916 570596 262922 570648
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 37918 565876 37924 565888
rect 3108 565848 37924 565876
rect 3108 565836 3114 565848
rect 37918 565836 37924 565848
rect 37976 565836 37982 565888
rect 403618 563048 403624 563100
rect 403676 563088 403682 563100
rect 580166 563088 580172 563100
rect 403676 563060 580172 563088
rect 403676 563048 403682 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 93486 559512 93492 559564
rect 93544 559552 93550 559564
rect 120718 559552 120724 559564
rect 93544 559524 120724 559552
rect 93544 559512 93550 559524
rect 120718 559512 120724 559524
rect 120776 559512 120782 559564
rect 193858 554752 193864 554804
rect 193916 554792 193922 554804
rect 196618 554792 196624 554804
rect 193916 554764 196624 554792
rect 193916 554752 193922 554764
rect 196618 554752 196624 554764
rect 196676 554752 196682 554804
rect 117958 553392 117964 553444
rect 118016 553432 118022 553444
rect 119338 553432 119344 553444
rect 118016 553404 119344 553432
rect 118016 553392 118022 553404
rect 119338 553392 119344 553404
rect 119396 553392 119402 553444
rect 90358 552508 90364 552560
rect 90416 552548 90422 552560
rect 93486 552548 93492 552560
rect 90416 552520 93492 552548
rect 90416 552508 90422 552520
rect 93486 552508 93492 552520
rect 93544 552508 93550 552560
rect 260190 552100 260196 552152
rect 260248 552140 260254 552152
rect 261478 552140 261484 552152
rect 260248 552112 261484 552140
rect 260248 552100 260254 552112
rect 261478 552100 261484 552112
rect 261536 552100 261542 552152
rect 258810 549992 258816 550044
rect 258868 550032 258874 550044
rect 260190 550032 260196 550044
rect 258868 550004 260196 550032
rect 258868 549992 258874 550004
rect 260190 549992 260196 550004
rect 260248 549992 260254 550044
rect 197998 545708 198004 545760
rect 198056 545748 198062 545760
rect 207658 545748 207664 545760
rect 198056 545720 207664 545748
rect 198056 545708 198062 545720
rect 207658 545708 207664 545720
rect 207716 545708 207722 545760
rect 256694 541968 256700 542020
rect 256752 542008 256758 542020
rect 258810 542008 258816 542020
rect 256752 541980 258816 542008
rect 256752 541968 256758 541980
rect 258810 541968 258816 541980
rect 258868 541968 258874 542020
rect 255958 538840 255964 538892
rect 256016 538880 256022 538892
rect 256694 538880 256700 538892
rect 256016 538852 256700 538880
rect 256016 538840 256022 538852
rect 256694 538840 256700 538852
rect 256752 538840 256758 538892
rect 116578 536800 116584 536852
rect 116636 536840 116642 536852
rect 117958 536840 117964 536852
rect 116636 536812 117964 536840
rect 116636 536800 116642 536812
rect 117958 536800 117964 536812
rect 118016 536800 118022 536852
rect 393958 536392 393964 536444
rect 394016 536432 394022 536444
rect 396626 536432 396632 536444
rect 394016 536404 396632 536432
rect 394016 536392 394022 536404
rect 396626 536392 396632 536404
rect 396684 536392 396690 536444
rect 115198 534080 115204 534132
rect 115256 534120 115262 534132
rect 116578 534120 116584 534132
rect 115256 534092 116584 534120
rect 115256 534080 115262 534092
rect 116578 534080 116584 534092
rect 116636 534080 116642 534132
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 6178 527184 6184 527196
rect 3016 527156 6184 527184
rect 3016 527144 3022 527156
rect 6178 527144 6184 527156
rect 6236 527144 6242 527196
rect 113818 525784 113824 525836
rect 113876 525824 113882 525836
rect 115198 525824 115204 525836
rect 113876 525796 115204 525824
rect 113876 525784 113882 525796
rect 115198 525784 115204 525796
rect 115256 525784 115262 525836
rect 181438 524464 181444 524476
rect 180766 524436 181444 524464
rect 177298 524356 177304 524408
rect 177356 524396 177362 524408
rect 180766 524396 180794 524436
rect 181438 524424 181444 524436
rect 181496 524424 181502 524476
rect 177356 524368 180794 524396
rect 177356 524356 177362 524368
rect 191098 520208 191104 520260
rect 191156 520248 191162 520260
rect 193858 520248 193864 520260
rect 191156 520220 193864 520248
rect 191156 520208 191162 520220
rect 193858 520208 193864 520220
rect 193916 520208 193922 520260
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 24118 514808 24124 514820
rect 3384 514780 24124 514808
rect 3384 514768 3390 514780
rect 24118 514768 24124 514780
rect 24176 514768 24182 514820
rect 253934 511776 253940 511828
rect 253992 511816 253998 511828
rect 255958 511816 255964 511828
rect 253992 511788 255964 511816
rect 253992 511776 253998 511788
rect 255958 511776 255964 511788
rect 256016 511776 256022 511828
rect 400858 510620 400864 510672
rect 400916 510660 400922 510672
rect 580166 510660 580172 510672
rect 400916 510632 580172 510660
rect 400916 510620 400922 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 251818 506472 251824 506524
rect 251876 506512 251882 506524
rect 253934 506512 253940 506524
rect 251876 506484 253940 506512
rect 251876 506472 251882 506484
rect 253934 506472 253940 506484
rect 253992 506472 253998 506524
rect 173158 505112 173164 505164
rect 173216 505152 173222 505164
rect 177298 505152 177304 505164
rect 173216 505124 177304 505152
rect 173216 505112 173222 505124
rect 177298 505112 177304 505124
rect 177356 505112 177362 505164
rect 195238 504364 195244 504416
rect 195296 504404 195302 504416
rect 197998 504404 198004 504416
rect 195296 504376 198004 504404
rect 195296 504364 195302 504376
rect 197998 504364 198004 504376
rect 198056 504364 198062 504416
rect 192478 490016 192484 490068
rect 192536 490056 192542 490068
rect 195238 490056 195244 490068
rect 192536 490028 195244 490056
rect 192536 490016 192542 490028
rect 195238 490016 195244 490028
rect 195296 490016 195302 490068
rect 112530 481652 112536 481704
rect 112588 481692 112594 481704
rect 113818 481692 113824 481704
rect 112588 481664 113824 481692
rect 112588 481652 112594 481664
rect 113818 481652 113824 481664
rect 113876 481652 113882 481704
rect 111058 476076 111064 476128
rect 111116 476116 111122 476128
rect 112530 476116 112536 476128
rect 111116 476088 112536 476116
rect 111116 476076 111122 476088
rect 112530 476076 112536 476088
rect 112588 476076 112594 476128
rect 171778 473016 171784 473068
rect 171836 473056 171842 473068
rect 173158 473056 173164 473068
rect 171836 473028 173164 473056
rect 171836 473016 171842 473028
rect 173158 473016 173164 473028
rect 173216 473016 173222 473068
rect 189074 470568 189080 470620
rect 189132 470608 189138 470620
rect 192478 470608 192484 470620
rect 189132 470580 192484 470608
rect 189132 470568 189138 470580
rect 192478 470568 192484 470580
rect 192536 470568 192542 470620
rect 182818 466420 182824 466472
rect 182876 466460 182882 466472
rect 189074 466460 189080 466472
rect 182876 466432 189080 466460
rect 182876 466420 182882 466432
rect 189074 466420 189080 466432
rect 189132 466420 189138 466472
rect 250162 466420 250168 466472
rect 250220 466460 250226 466472
rect 251818 466460 251824 466472
rect 250220 466432 251824 466460
rect 250220 466420 250226 466432
rect 251818 466420 251824 466432
rect 251876 466420 251882 466472
rect 248414 462952 248420 463004
rect 248472 462992 248478 463004
rect 250162 462992 250168 463004
rect 248472 462964 250168 462992
rect 248472 462952 248478 462964
rect 250162 462952 250168 462964
rect 250220 462952 250226 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4982 462584 4988 462596
rect 2832 462556 4988 462584
rect 2832 462544 2838 462556
rect 4982 462544 4988 462556
rect 5040 462544 5046 462596
rect 109678 459552 109684 459604
rect 109736 459592 109742 459604
rect 111058 459592 111064 459604
rect 109736 459564 111064 459592
rect 109736 459552 109742 459564
rect 111058 459552 111064 459564
rect 111116 459552 111122 459604
rect 179414 459552 179420 459604
rect 179472 459592 179478 459604
rect 182818 459592 182824 459604
rect 179472 459564 182824 459592
rect 179472 459552 179478 459564
rect 182818 459552 182824 459564
rect 182876 459552 182882 459604
rect 245746 459552 245752 459604
rect 245804 459592 245810 459604
rect 248414 459592 248420 459604
rect 245804 459564 248420 459592
rect 245804 459552 245810 459564
rect 248414 459552 248420 459564
rect 248472 459552 248478 459604
rect 399478 456764 399484 456816
rect 399536 456804 399542 456816
rect 579982 456804 579988 456816
rect 399536 456776 579988 456804
rect 399536 456764 399542 456776
rect 579982 456764 579988 456776
rect 580040 456764 580046 456816
rect 244918 455404 244924 455456
rect 244976 455444 244982 455456
rect 245746 455444 245752 455456
rect 244976 455416 245752 455444
rect 244976 455404 244982 455416
rect 245746 455404 245752 455416
rect 245804 455404 245810 455456
rect 177298 452548 177304 452600
rect 177356 452588 177362 452600
rect 179414 452588 179420 452600
rect 177356 452560 179420 452588
rect 177356 452548 177362 452560
rect 179414 452548 179420 452560
rect 179472 452548 179478 452600
rect 84194 452072 84200 452124
rect 84252 452112 84258 452124
rect 90358 452112 90364 452124
rect 84252 452084 90364 452112
rect 84252 452072 84258 452084
rect 90358 452072 90364 452084
rect 90416 452072 90422 452124
rect 75178 447788 75184 447840
rect 75236 447828 75242 447840
rect 84194 447828 84200 447840
rect 75236 447800 84200 447828
rect 75236 447788 75242 447800
rect 84194 447788 84200 447800
rect 84252 447788 84258 447840
rect 170398 447040 170404 447092
rect 170456 447080 170462 447092
rect 171778 447080 171784 447092
rect 170456 447052 171784 447080
rect 170456 447040 170462 447052
rect 171778 447040 171784 447052
rect 171836 447040 171842 447092
rect 170398 437492 170404 437504
rect 168392 437464 170404 437492
rect 166994 437384 167000 437436
rect 167052 437424 167058 437436
rect 168392 437424 168420 437464
rect 170398 437452 170404 437464
rect 170456 437452 170462 437504
rect 167052 437396 168420 437424
rect 167052 437384 167058 437396
rect 151078 436704 151084 436756
rect 151136 436744 151142 436756
rect 177298 436744 177304 436756
rect 151136 436716 177304 436744
rect 151136 436704 151142 436716
rect 177298 436704 177304 436716
rect 177356 436704 177362 436756
rect 166902 433344 166908 433356
rect 164252 433316 166908 433344
rect 163590 433236 163596 433288
rect 163648 433276 163654 433288
rect 164252 433276 164280 433316
rect 166902 433304 166908 433316
rect 166960 433304 166966 433356
rect 163648 433248 164280 433276
rect 163648 433236 163654 433248
rect 134702 431196 134708 431248
rect 134760 431236 134766 431248
rect 151078 431236 151084 431248
rect 134760 431208 151084 431236
rect 134760 431196 134766 431208
rect 151078 431196 151084 431208
rect 151136 431196 151142 431248
rect 107654 430584 107660 430636
rect 107712 430624 107718 430636
rect 109678 430624 109684 430636
rect 107712 430596 109684 430624
rect 107712 430584 107718 430596
rect 109678 430584 109684 430596
rect 109736 430584 109742 430636
rect 171502 429836 171508 429888
rect 171560 429876 171566 429888
rect 191098 429876 191104 429888
rect 171560 429848 191104 429876
rect 171560 429836 171566 429848
rect 191098 429836 191104 429848
rect 191156 429836 191162 429888
rect 106182 427116 106188 427168
rect 106240 427156 106246 427168
rect 107654 427156 107660 427168
rect 106240 427128 107660 427156
rect 106240 427116 106246 427128
rect 107654 427116 107660 427128
rect 107712 427116 107718 427168
rect 163498 425688 163504 425740
rect 163556 425728 163562 425740
rect 171502 425728 171508 425740
rect 163556 425700 171508 425728
rect 163556 425688 163562 425700
rect 171502 425688 171508 425700
rect 171560 425688 171566 425740
rect 103514 423240 103520 423292
rect 103572 423280 103578 423292
rect 106182 423280 106188 423292
rect 103572 423252 106188 423280
rect 103572 423240 103578 423252
rect 106182 423240 106188 423252
rect 106240 423240 106246 423292
rect 131758 422288 131764 422340
rect 131816 422328 131822 422340
rect 134702 422328 134708 422340
rect 131816 422300 134708 422328
rect 131816 422288 131822 422300
rect 134702 422288 134708 422300
rect 134760 422288 134766 422340
rect 398098 418140 398104 418192
rect 398156 418180 398162 418192
rect 580074 418180 580080 418192
rect 398156 418152 580080 418180
rect 398156 418140 398162 418152
rect 580074 418140 580080 418152
rect 580132 418140 580138 418192
rect 101398 417664 101404 417716
rect 101456 417704 101462 417716
rect 103514 417704 103520 417716
rect 101456 417676 103520 417704
rect 101456 417664 101462 417676
rect 103514 417664 103520 417676
rect 103572 417664 103578 417716
rect 243538 416712 243544 416764
rect 243596 416752 243602 416764
rect 244918 416752 244924 416764
rect 243596 416724 244924 416752
rect 243596 416712 243602 416724
rect 244918 416712 244924 416724
rect 244976 416712 244982 416764
rect 160738 413992 160744 414044
rect 160796 414032 160802 414044
rect 163590 414032 163596 414044
rect 160796 414004 163596 414032
rect 160796 413992 160802 414004
rect 163590 413992 163596 414004
rect 163648 413992 163654 414044
rect 113174 413244 113180 413296
rect 113232 413284 113238 413296
rect 131758 413284 131764 413296
rect 113232 413256 131764 413284
rect 113232 413244 113238 413256
rect 131758 413244 131764 413256
rect 131816 413244 131822 413296
rect 3234 410456 3240 410508
rect 3292 410496 3298 410508
rect 8938 410496 8944 410508
rect 3292 410468 8944 410496
rect 3292 410456 3298 410468
rect 8938 410456 8944 410468
rect 8996 410456 9002 410508
rect 95326 407736 95332 407788
rect 95384 407776 95390 407788
rect 113174 407776 113180 407788
rect 95384 407748 113180 407776
rect 95384 407736 95390 407748
rect 113174 407736 113180 407748
rect 113232 407736 113238 407788
rect 160830 407056 160836 407108
rect 160888 407096 160894 407108
rect 163498 407096 163504 407108
rect 160888 407068 163504 407096
rect 160888 407056 160894 407068
rect 163498 407056 163504 407068
rect 163556 407056 163562 407108
rect 101398 405736 101404 405748
rect 98012 405708 101404 405736
rect 97442 405628 97448 405680
rect 97500 405668 97506 405680
rect 98012 405668 98040 405708
rect 101398 405696 101404 405708
rect 101456 405696 101462 405748
rect 97500 405640 98040 405668
rect 97500 405628 97506 405640
rect 418798 404336 418804 404388
rect 418856 404376 418862 404388
rect 580074 404376 580080 404388
rect 418856 404348 580080 404376
rect 418856 404336 418862 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 75270 403588 75276 403640
rect 75328 403628 75334 403640
rect 95326 403628 95332 403640
rect 75328 403600 95332 403628
rect 75328 403588 75334 403600
rect 95326 403588 95332 403600
rect 95384 403588 95390 403640
rect 236638 403588 236644 403640
rect 236696 403628 236702 403640
rect 243538 403628 243544 403640
rect 236696 403600 243544 403628
rect 236696 403588 236702 403600
rect 243538 403588 243544 403600
rect 243596 403588 243602 403640
rect 148318 402228 148324 402280
rect 148376 402268 148382 402280
rect 160830 402268 160836 402280
rect 148376 402240 160836 402268
rect 148376 402228 148382 402240
rect 160830 402228 160836 402240
rect 160888 402228 160894 402280
rect 96062 401616 96068 401668
rect 96120 401656 96126 401668
rect 97442 401656 97448 401668
rect 96120 401628 97448 401656
rect 96120 401616 96126 401628
rect 97442 401616 97448 401628
rect 97500 401616 97506 401668
rect 94498 397808 94504 397860
rect 94556 397848 94562 397860
rect 96062 397848 96068 397860
rect 94556 397820 96068 397848
rect 94556 397808 94562 397820
rect 96062 397808 96068 397820
rect 96120 397808 96126 397860
rect 69658 396720 69664 396772
rect 69716 396760 69722 396772
rect 136634 396760 136640 396772
rect 69716 396732 136640 396760
rect 69716 396720 69722 396732
rect 136634 396720 136640 396732
rect 136692 396720 136698 396772
rect 233878 395972 233884 396024
rect 233936 396012 233942 396024
rect 236638 396012 236644 396024
rect 233936 395984 236644 396012
rect 233936 395972 233942 395984
rect 236638 395972 236644 395984
rect 236696 395972 236702 396024
rect 72418 391960 72424 392012
rect 72476 392000 72482 392012
rect 75178 392000 75184 392012
rect 72476 391972 75184 392000
rect 72476 391960 72482 391972
rect 75178 391960 75184 391972
rect 75236 391960 75242 392012
rect 92474 390736 92480 390788
rect 92532 390776 92538 390788
rect 94498 390776 94504 390788
rect 92532 390748 94504 390776
rect 92532 390736 92538 390748
rect 94498 390736 94504 390748
rect 94556 390736 94562 390788
rect 90082 385704 90088 385756
rect 90140 385744 90146 385756
rect 92474 385744 92480 385756
rect 90140 385716 92480 385744
rect 90140 385704 90146 385716
rect 92474 385704 92480 385716
rect 92532 385704 92538 385756
rect 68278 384956 68284 385008
rect 68336 384996 68342 385008
rect 69658 384996 69664 385008
rect 68336 384968 69664 384996
rect 68336 384956 68342 384968
rect 69658 384956 69664 384968
rect 69716 384956 69722 385008
rect 86218 382236 86224 382288
rect 86276 382276 86282 382288
rect 90082 382276 90088 382288
rect 86276 382248 90088 382276
rect 86276 382236 86282 382248
rect 90082 382236 90088 382248
rect 90140 382236 90146 382288
rect 396810 378156 396816 378208
rect 396868 378196 396874 378208
rect 580074 378196 580080 378208
rect 396868 378168 580080 378196
rect 396868 378156 396874 378168
rect 580074 378156 580080 378168
rect 580132 378156 580138 378208
rect 3234 371220 3240 371272
rect 3292 371260 3298 371272
rect 10410 371260 10416 371272
rect 3292 371232 10416 371260
rect 3292 371220 3298 371232
rect 10410 371220 10416 371232
rect 10468 371220 10474 371272
rect 59262 370472 59268 370524
rect 59320 370512 59326 370524
rect 72418 370512 72424 370524
rect 59320 370484 72424 370512
rect 59320 370472 59326 370484
rect 72418 370472 72424 370484
rect 72476 370472 72482 370524
rect 159358 366732 159364 366784
rect 159416 366772 159422 366784
rect 160738 366772 160744 366784
rect 159416 366744 160744 366772
rect 159416 366732 159422 366744
rect 160738 366732 160744 366744
rect 160796 366732 160802 366784
rect 46934 366324 46940 366376
rect 46992 366364 46998 366376
rect 59262 366364 59268 366376
rect 46992 366336 59268 366364
rect 46992 366324 46998 366336
rect 59262 366324 59268 366336
rect 59320 366324 59326 366376
rect 398190 364352 398196 364404
rect 398248 364392 398254 364404
rect 579798 364392 579804 364404
rect 398248 364364 579804 364392
rect 398248 364352 398254 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 45094 360952 45100 361004
rect 45152 360992 45158 361004
rect 46934 360992 46940 361004
rect 45152 360964 46940 360992
rect 45152 360952 45158 360964
rect 46934 360952 46940 360964
rect 46992 360952 46998 361004
rect 84838 358980 84844 359032
rect 84896 359020 84902 359032
rect 86218 359020 86224 359032
rect 84896 358992 86224 359020
rect 84896 358980 84902 358992
rect 86218 358980 86224 358992
rect 86276 358980 86282 359032
rect 65426 358776 65432 358828
rect 65484 358816 65490 358828
rect 68278 358816 68284 358828
rect 65484 358788 68284 358816
rect 65484 358776 65490 358788
rect 68278 358776 68284 358788
rect 68336 358776 68342 358828
rect 64138 358096 64144 358148
rect 64196 358136 64202 358148
rect 65426 358136 65432 358148
rect 64196 358108 65432 358136
rect 64196 358096 64202 358108
rect 65426 358096 65432 358108
rect 65484 358096 65490 358148
rect 3234 357416 3240 357468
rect 3292 357456 3298 357468
rect 22738 357456 22744 357468
rect 3292 357428 22744 357456
rect 3292 357416 3298 357428
rect 22738 357416 22744 357428
rect 22796 357416 22802 357468
rect 157978 355988 157984 356040
rect 158036 356028 158042 356040
rect 159358 356028 159364 356040
rect 158036 356000 159364 356028
rect 158036 355988 158042 356000
rect 159358 355988 159364 356000
rect 159416 355988 159422 356040
rect 71866 353268 71872 353320
rect 71924 353308 71930 353320
rect 75270 353308 75276 353320
rect 71924 353280 75276 353308
rect 71924 353268 71930 353280
rect 75270 353268 75276 353280
rect 75328 353268 75334 353320
rect 145558 353268 145564 353320
rect 145616 353308 145622 353320
rect 148318 353308 148324 353320
rect 145616 353280 148324 353308
rect 145616 353268 145622 353280
rect 148318 353268 148324 353280
rect 148376 353268 148382 353320
rect 84838 351948 84844 351960
rect 84166 351920 84844 351948
rect 82354 351840 82360 351892
rect 82412 351880 82418 351892
rect 84166 351880 84194 351920
rect 84838 351908 84844 351920
rect 84896 351908 84902 351960
rect 417418 351908 417424 351960
rect 417476 351948 417482 351960
rect 580074 351948 580080 351960
rect 417476 351920 580080 351948
rect 417476 351908 417482 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 82412 351852 84194 351880
rect 82412 351840 82418 351852
rect 228358 349800 228364 349852
rect 228416 349840 228422 349852
rect 233878 349840 233884 349852
rect 228416 349812 233884 349840
rect 228416 349800 228422 349812
rect 233878 349800 233884 349812
rect 233936 349800 233942 349852
rect 80698 349120 80704 349172
rect 80756 349160 80762 349172
rect 82354 349160 82360 349172
rect 80756 349132 82360 349160
rect 80756 349120 80762 349132
rect 82354 349120 82360 349132
rect 82412 349120 82418 349172
rect 63862 345652 63868 345704
rect 63920 345692 63926 345704
rect 71866 345692 71872 345704
rect 63920 345664 71872 345692
rect 63920 345652 63926 345664
rect 71866 345652 71872 345664
rect 71924 345652 71930 345704
rect 61378 339192 61384 339244
rect 61436 339232 61442 339244
rect 63862 339232 63868 339244
rect 61436 339204 63868 339232
rect 61436 339192 61442 339204
rect 63862 339192 63868 339204
rect 63920 339192 63926 339244
rect 225598 338036 225604 338088
rect 225656 338076 225662 338088
rect 228358 338076 228364 338088
rect 225656 338048 228364 338076
rect 225656 338036 225662 338048
rect 228358 338036 228364 338048
rect 228416 338036 228422 338088
rect 140406 337356 140412 337408
rect 140464 337396 140470 337408
rect 145558 337396 145564 337408
rect 140464 337368 145564 337396
rect 140464 337356 140470 337368
rect 145558 337356 145564 337368
rect 145616 337356 145622 337408
rect 156690 332596 156696 332648
rect 156748 332636 156754 332648
rect 157978 332636 157984 332648
rect 156748 332608 157984 332636
rect 156748 332596 156754 332608
rect 157978 332596 157984 332608
rect 158036 332596 158042 332648
rect 62850 331848 62856 331900
rect 62908 331888 62914 331900
rect 88334 331888 88340 331900
rect 62908 331860 88340 331888
rect 62908 331848 62914 331860
rect 88334 331848 88340 331860
rect 88392 331848 88398 331900
rect 135898 328856 135904 328908
rect 135956 328896 135962 328908
rect 140406 328896 140412 328908
rect 135956 328868 140412 328896
rect 135956 328856 135962 328868
rect 140406 328856 140412 328868
rect 140464 328856 140470 328908
rect 155218 328040 155224 328092
rect 155276 328080 155282 328092
rect 156690 328080 156696 328092
rect 155276 328052 156696 328080
rect 155276 328040 155282 328052
rect 156690 328040 156696 328052
rect 156748 328040 156754 328092
rect 396994 324300 397000 324352
rect 397052 324340 397058 324352
rect 580074 324340 580080 324352
rect 397052 324312 580080 324340
rect 397052 324300 397058 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 79502 320152 79508 320204
rect 79560 320192 79566 320204
rect 80698 320192 80704 320204
rect 79560 320164 80704 320192
rect 79560 320152 79566 320164
rect 80698 320152 80704 320164
rect 80756 320152 80762 320204
rect 62758 319404 62764 319456
rect 62816 319444 62822 319456
rect 64138 319444 64144 319456
rect 62816 319416 64144 319444
rect 62816 319404 62822 319416
rect 64138 319404 64144 319416
rect 64196 319404 64202 319456
rect 3234 318792 3240 318844
rect 3292 318832 3298 318844
rect 33778 318832 33784 318844
rect 3292 318804 33784 318832
rect 3292 318792 3298 318804
rect 33778 318792 33784 318804
rect 33836 318792 33842 318844
rect 153838 318724 153844 318776
rect 153896 318764 153902 318776
rect 155218 318764 155224 318776
rect 153896 318736 155224 318764
rect 153896 318724 153902 318736
rect 155218 318724 155224 318736
rect 155276 318724 155282 318776
rect 61470 318384 61476 318436
rect 61528 318424 61534 318436
rect 62850 318424 62856 318436
rect 61528 318396 62856 318424
rect 61528 318384 61534 318396
rect 62850 318384 62856 318396
rect 62908 318384 62914 318436
rect 78122 318316 78128 318368
rect 78180 318356 78186 318368
rect 79502 318356 79508 318368
rect 78180 318328 79508 318356
rect 78180 318316 78186 318328
rect 79502 318316 79508 318328
rect 79560 318316 79566 318368
rect 224218 317364 224224 317416
rect 224276 317404 224282 317416
rect 225598 317404 225604 317416
rect 224276 317376 225604 317404
rect 224276 317364 224282 317376
rect 225598 317364 225604 317376
rect 225656 317364 225662 317416
rect 73154 315256 73160 315308
rect 73212 315296 73218 315308
rect 78122 315296 78128 315308
rect 73212 315268 78128 315296
rect 73212 315256 73218 315268
rect 78122 315256 78128 315268
rect 78180 315256 78186 315308
rect 84838 315256 84844 315308
rect 84896 315296 84902 315308
rect 104894 315296 104900 315308
rect 84896 315268 104900 315296
rect 84896 315256 84902 315268
rect 104894 315256 104900 315268
rect 104952 315256 104958 315308
rect 58618 314644 58624 314696
rect 58676 314684 58682 314696
rect 61378 314684 61384 314696
rect 58676 314656 61384 314684
rect 58676 314644 58682 314656
rect 61378 314644 61384 314656
rect 61436 314644 61442 314696
rect 71038 313284 71044 313336
rect 71096 313324 71102 313336
rect 73154 313324 73160 313336
rect 71096 313296 73160 313324
rect 71096 313284 71102 313296
rect 73154 313284 73160 313296
rect 73212 313284 73218 313336
rect 398282 311856 398288 311908
rect 398340 311896 398346 311908
rect 580074 311896 580080 311908
rect 398340 311868 580080 311896
rect 398340 311856 398346 311868
rect 580074 311856 580080 311868
rect 580132 311856 580138 311908
rect 59998 311176 60004 311228
rect 60056 311216 60062 311228
rect 61470 311216 61476 311228
rect 60056 311188 61476 311216
rect 60056 311176 60062 311188
rect 61470 311176 61476 311188
rect 61528 311176 61534 311228
rect 102778 308388 102784 308440
rect 102836 308428 102842 308440
rect 135898 308428 135904 308440
rect 102836 308400 135904 308428
rect 102836 308388 102842 308400
rect 135898 308388 135904 308400
rect 135956 308388 135962 308440
rect 153838 307816 153844 307828
rect 151786 307788 153844 307816
rect 151078 307708 151084 307760
rect 151136 307748 151142 307760
rect 151786 307748 151814 307788
rect 153838 307776 153844 307788
rect 153896 307776 153902 307828
rect 151136 307720 151814 307748
rect 151136 307708 151142 307720
rect 69658 304988 69664 305040
rect 69716 305028 69722 305040
rect 71038 305028 71044 305040
rect 69716 305000 71044 305028
rect 69716 304988 69722 305000
rect 71038 304988 71044 305000
rect 71096 304988 71102 305040
rect 224218 303668 224224 303680
rect 222212 303640 224224 303668
rect 220814 303560 220820 303612
rect 220872 303600 220878 303612
rect 222212 303600 222240 303640
rect 224218 303628 224224 303640
rect 224276 303628 224282 303680
rect 220872 303572 222240 303600
rect 220872 303560 220878 303572
rect 68278 302200 68284 302252
rect 68336 302240 68342 302252
rect 69658 302240 69664 302252
rect 68336 302212 69664 302240
rect 68336 302200 68342 302212
rect 69658 302200 69664 302212
rect 69716 302200 69722 302252
rect 220078 301112 220084 301164
rect 220136 301152 220142 301164
rect 220814 301152 220820 301164
rect 220136 301124 220820 301152
rect 220136 301112 220142 301124
rect 220814 301112 220820 301124
rect 220872 301112 220878 301164
rect 60826 299412 60832 299464
rect 60884 299452 60890 299464
rect 62758 299452 62764 299464
rect 60884 299424 62764 299452
rect 60884 299412 60890 299424
rect 62758 299412 62764 299424
rect 62816 299412 62822 299464
rect 414658 298120 414664 298172
rect 414716 298160 414722 298172
rect 580074 298160 580080 298172
rect 414716 298132 580080 298160
rect 414716 298120 414722 298132
rect 580074 298120 580080 298132
rect 580132 298120 580138 298172
rect 97718 297372 97724 297424
rect 97776 297412 97782 297424
rect 102778 297412 102784 297424
rect 97776 297384 102784 297412
rect 97776 297372 97782 297384
rect 102778 297372 102784 297384
rect 102836 297372 102842 297424
rect 87598 294584 87604 294636
rect 87656 294624 87662 294636
rect 97718 294624 97724 294636
rect 87656 294596 97724 294624
rect 87656 294584 87662 294596
rect 97718 294584 97724 294596
rect 97776 294584 97782 294636
rect 66254 294176 66260 294228
rect 66312 294216 66318 294228
rect 68278 294216 68284 294228
rect 66312 294188 68284 294216
rect 66312 294176 66318 294188
rect 68278 294176 68284 294188
rect 68336 294176 68342 294228
rect 60090 293972 60096 294024
rect 60148 294012 60154 294024
rect 60826 294012 60832 294024
rect 60148 293984 60832 294012
rect 60148 293972 60154 293984
rect 60826 293972 60832 293984
rect 60884 293972 60890 294024
rect 2774 292612 2780 292664
rect 2832 292652 2838 292664
rect 5074 292652 5080 292664
rect 2832 292624 5080 292652
rect 2832 292612 2838 292624
rect 5074 292612 5080 292624
rect 5132 292612 5138 292664
rect 63494 292612 63500 292664
rect 63552 292652 63558 292664
rect 66254 292652 66260 292664
rect 63552 292624 66260 292652
rect 63552 292612 63558 292624
rect 66254 292612 66260 292624
rect 66312 292612 66318 292664
rect 53834 291796 53840 291848
rect 53892 291836 53898 291848
rect 63494 291836 63500 291848
rect 53892 291808 63500 291836
rect 53892 291796 53898 291808
rect 63494 291796 63500 291808
rect 63552 291796 63558 291848
rect 220078 291224 220084 291236
rect 213932 291196 220084 291224
rect 213822 291116 213828 291168
rect 213880 291156 213886 291168
rect 213932 291156 213960 291196
rect 220078 291184 220084 291196
rect 220136 291184 220142 291236
rect 213880 291128 213960 291156
rect 213880 291116 213886 291128
rect 58710 290368 58716 290420
rect 58768 290408 58774 290420
rect 59998 290408 60004 290420
rect 58768 290380 60004 290408
rect 58768 290368 58774 290380
rect 59998 290368 60004 290380
rect 60056 290368 60062 290420
rect 53834 289864 53840 289876
rect 52472 289836 53840 289864
rect 51810 289756 51816 289808
rect 51868 289796 51874 289808
rect 52472 289796 52500 289836
rect 53834 289824 53840 289836
rect 53892 289824 53898 289876
rect 51868 289768 52500 289796
rect 51868 289756 51874 289768
rect 211154 288872 211160 288924
rect 211212 288912 211218 288924
rect 213822 288912 213828 288924
rect 211212 288884 213828 288912
rect 211212 288872 211218 288884
rect 213822 288872 213828 288884
rect 213880 288872 213886 288924
rect 57238 287648 57244 287700
rect 57296 287688 57302 287700
rect 71774 287688 71780 287700
rect 57296 287660 71780 287688
rect 57296 287648 57302 287660
rect 71774 287648 71780 287660
rect 71832 287648 71838 287700
rect 82814 284928 82820 284980
rect 82872 284968 82878 284980
rect 87598 284968 87604 284980
rect 82872 284940 87604 284968
rect 82872 284928 82878 284940
rect 87598 284928 87604 284940
rect 87656 284928 87662 284980
rect 58710 284356 58716 284368
rect 56612 284328 58716 284356
rect 55582 284248 55588 284300
rect 55640 284288 55646 284300
rect 56612 284288 56640 284328
rect 58710 284316 58716 284328
rect 58768 284316 58774 284368
rect 84838 284356 84844 284368
rect 84166 284328 84844 284356
rect 55640 284260 56640 284288
rect 55640 284248 55646 284260
rect 82078 284248 82084 284300
rect 82136 284288 82142 284300
rect 84166 284288 84194 284328
rect 84838 284316 84844 284328
rect 84896 284316 84902 284368
rect 82136 284260 84194 284288
rect 82136 284248 82142 284260
rect 207014 283976 207020 284028
rect 207072 284016 207078 284028
rect 211154 284016 211160 284028
rect 207072 283988 211160 284016
rect 207072 283976 207078 283988
rect 211154 283976 211160 283988
rect 211212 283976 211218 284028
rect 57974 282888 57980 282940
rect 58032 282928 58038 282940
rect 60090 282928 60096 282940
rect 58032 282900 60096 282928
rect 58032 282888 58038 282900
rect 60090 282888 60096 282900
rect 60148 282888 60154 282940
rect 66898 282140 66904 282192
rect 66956 282180 66962 282192
rect 82814 282180 82820 282192
rect 66956 282152 82820 282180
rect 66956 282140 66962 282152
rect 82814 282140 82820 282152
rect 82872 282140 82878 282192
rect 148318 281256 148324 281308
rect 148376 281296 148382 281308
rect 151078 281296 151084 281308
rect 148376 281268 151084 281296
rect 148376 281256 148382 281268
rect 151078 281256 151084 281268
rect 151136 281256 151142 281308
rect 54202 281120 54208 281172
rect 54260 281160 54266 281172
rect 55582 281160 55588 281172
rect 54260 281132 55588 281160
rect 54260 281120 54266 281132
rect 55582 281120 55588 281132
rect 55640 281120 55646 281172
rect 53282 280780 53288 280832
rect 53340 280820 53346 280832
rect 169754 280820 169760 280832
rect 53340 280792 169760 280820
rect 53340 280780 53346 280792
rect 169754 280780 169760 280792
rect 169812 280780 169818 280832
rect 49694 280168 49700 280220
rect 49752 280208 49758 280220
rect 51810 280208 51816 280220
rect 49752 280180 51816 280208
rect 49752 280168 49758 280180
rect 51810 280168 51816 280180
rect 51868 280168 51874 280220
rect 53098 278808 53104 278860
rect 53156 278848 53162 278860
rect 54202 278848 54208 278860
rect 53156 278820 54208 278848
rect 53156 278808 53162 278820
rect 54202 278808 54208 278820
rect 54260 278808 54266 278860
rect 54478 278740 54484 278792
rect 54536 278780 54542 278792
rect 57882 278780 57888 278792
rect 54536 278752 57888 278780
rect 54536 278740 54542 278752
rect 57882 278740 57888 278752
rect 57940 278740 57946 278792
rect 204162 278264 204168 278316
rect 204220 278304 204226 278316
rect 207014 278304 207020 278316
rect 204220 278276 207020 278304
rect 204220 278264 204226 278276
rect 207014 278264 207020 278276
rect 207072 278264 207078 278316
rect 48958 278128 48964 278180
rect 49016 278168 49022 278180
rect 49694 278168 49700 278180
rect 49016 278140 49700 278168
rect 49016 278128 49022 278140
rect 49694 278128 49700 278140
rect 49752 278128 49758 278180
rect 46934 277992 46940 278044
rect 46992 278032 46998 278044
rect 58618 278032 58624 278044
rect 46992 278004 58624 278032
rect 46992 277992 46998 278004
rect 58618 277992 58624 278004
rect 58676 277992 58682 278044
rect 57238 277420 57244 277432
rect 55232 277392 57244 277420
rect 53834 277312 53840 277364
rect 53892 277352 53898 277364
rect 55232 277352 55260 277392
rect 57238 277380 57244 277392
rect 57296 277380 57302 277432
rect 53892 277324 55260 277352
rect 53892 277312 53898 277324
rect 55858 276632 55864 276684
rect 55916 276672 55922 276684
rect 82078 276672 82084 276684
rect 55916 276644 82084 276672
rect 55916 276632 55922 276644
rect 82078 276632 82084 276644
rect 82136 276632 82142 276684
rect 63494 275068 63500 275120
rect 63552 275108 63558 275120
rect 66898 275108 66904 275120
rect 63552 275080 66904 275108
rect 63552 275068 63558 275080
rect 66898 275068 66904 275080
rect 66956 275068 66962 275120
rect 44910 274660 44916 274712
rect 44968 274700 44974 274712
rect 46934 274700 46940 274712
rect 44968 274672 46940 274700
rect 44968 274660 44974 274672
rect 46934 274660 46940 274672
rect 46992 274660 46998 274712
rect 53190 274660 53196 274712
rect 53248 274700 53254 274712
rect 53834 274700 53840 274712
rect 53248 274672 53840 274700
rect 53248 274660 53254 274672
rect 53834 274660 53840 274672
rect 53892 274660 53898 274712
rect 201494 274660 201500 274712
rect 201552 274700 201558 274712
rect 204162 274700 204168 274712
rect 201552 274672 204168 274700
rect 201552 274660 201558 274672
rect 204162 274660 204168 274672
rect 204220 274660 204226 274712
rect 51718 272008 51724 272060
rect 51776 272048 51782 272060
rect 53098 272048 53104 272060
rect 51776 272020 53104 272048
rect 51776 272008 51782 272020
rect 53098 272008 53104 272020
rect 53156 272008 53162 272060
rect 504358 271872 504364 271924
rect 504416 271912 504422 271924
rect 579798 271912 579804 271924
rect 504416 271884 579804 271912
rect 504416 271872 504422 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 200758 270920 200764 270972
rect 200816 270960 200822 270972
rect 201494 270960 201500 270972
rect 200816 270932 201500 270960
rect 200816 270920 200822 270932
rect 201494 270920 201500 270932
rect 201552 270920 201558 270972
rect 51074 270444 51080 270496
rect 51132 270484 51138 270496
rect 53282 270484 53288 270496
rect 51132 270456 53288 270484
rect 51132 270444 51138 270456
rect 53282 270444 53288 270456
rect 53340 270444 53346 270496
rect 60550 268608 60556 268660
rect 60608 268648 60614 268660
rect 63494 268648 63500 268660
rect 60608 268620 63500 268648
rect 60608 268608 60614 268620
rect 63494 268608 63500 268620
rect 63552 268608 63558 268660
rect 53190 266432 53196 266484
rect 53248 266472 53254 266484
rect 54478 266472 54484 266484
rect 53248 266444 54484 266472
rect 53248 266432 53254 266444
rect 54478 266432 54484 266444
rect 54536 266432 54542 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 20070 266404 20076 266416
rect 3108 266376 20076 266404
rect 3108 266364 3114 266376
rect 20070 266364 20076 266376
rect 20128 266364 20134 266416
rect 51074 266404 51080 266416
rect 49712 266376 51080 266404
rect 48314 266296 48320 266348
rect 48372 266336 48378 266348
rect 49712 266336 49740 266376
rect 51074 266364 51080 266376
rect 51132 266364 51138 266416
rect 54202 266364 54208 266416
rect 54260 266404 54266 266416
rect 55858 266404 55864 266416
rect 54260 266376 55864 266404
rect 54260 266364 54266 266376
rect 55858 266364 55864 266376
rect 55916 266364 55922 266416
rect 197998 266364 198004 266416
rect 198056 266404 198062 266416
rect 200758 266404 200764 266416
rect 198056 266376 200764 266404
rect 198056 266364 198062 266376
rect 200758 266364 200764 266376
rect 200816 266364 200822 266416
rect 48372 266308 49740 266336
rect 48372 266296 48378 266308
rect 49694 263576 49700 263628
rect 49752 263616 49758 263628
rect 51718 263616 51724 263628
rect 49752 263588 51724 263616
rect 49752 263576 49758 263588
rect 51718 263576 51724 263588
rect 51776 263576 51782 263628
rect 53282 263576 53288 263628
rect 53340 263616 53346 263628
rect 54202 263616 54208 263628
rect 53340 263588 54208 263616
rect 53340 263576 53346 263588
rect 54202 263576 54208 263588
rect 54260 263576 54266 263628
rect 146938 262896 146944 262948
rect 146996 262936 147002 262948
rect 148318 262936 148324 262948
rect 146996 262908 148324 262936
rect 146996 262896 147002 262908
rect 148318 262896 148324 262908
rect 148376 262896 148382 262948
rect 53374 262828 53380 262880
rect 53432 262868 53438 262880
rect 60550 262868 60556 262880
rect 53432 262840 60556 262868
rect 53432 262828 53438 262840
rect 60550 262828 60556 262840
rect 60608 262828 60614 262880
rect 45738 259224 45744 259276
rect 45796 259264 45802 259276
rect 48222 259264 48228 259276
rect 45796 259236 48228 259264
rect 45796 259224 45802 259236
rect 48222 259224 48228 259236
rect 48280 259224 48286 259276
rect 46934 258544 46940 258596
rect 46992 258584 46998 258596
rect 49694 258584 49700 258596
rect 46992 258556 49700 258584
rect 46992 258544 46998 258556
rect 49694 258544 49700 258556
rect 49752 258544 49758 258596
rect 398374 258068 398380 258120
rect 398432 258108 398438 258120
rect 579982 258108 579988 258120
rect 398432 258080 579988 258108
rect 398432 258068 398438 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 48222 256776 48228 256828
rect 48280 256816 48286 256828
rect 53374 256816 53380 256828
rect 48280 256788 53380 256816
rect 48280 256776 48286 256788
rect 53374 256776 53380 256788
rect 53432 256776 53438 256828
rect 53282 256748 53288 256760
rect 51092 256720 53288 256748
rect 50430 256640 50436 256692
rect 50488 256680 50494 256692
rect 51092 256680 51120 256720
rect 53282 256708 53288 256720
rect 53340 256708 53346 256760
rect 50488 256652 51120 256680
rect 50488 256640 50494 256652
rect 45554 255280 45560 255332
rect 45612 255320 45618 255332
rect 46934 255320 46940 255332
rect 45612 255292 46940 255320
rect 45612 255280 45618 255292
rect 46934 255280 46940 255292
rect 46992 255280 46998 255332
rect 45002 254260 45008 254312
rect 45060 254300 45066 254312
rect 48222 254300 48228 254312
rect 45060 254272 48228 254300
rect 45060 254260 45066 254272
rect 48222 254260 48228 254272
rect 48280 254260 48286 254312
rect 47578 253988 47584 254040
rect 47636 254028 47642 254040
rect 50430 254028 50436 254040
rect 47636 254000 50436 254028
rect 47636 253988 47642 254000
rect 50430 253988 50436 254000
rect 50488 253988 50494 254040
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 22830 253960 22836 253972
rect 3200 253932 22836 253960
rect 3200 253920 3206 253932
rect 22830 253920 22836 253932
rect 22888 253920 22894 253972
rect 46934 253920 46940 253972
rect 46992 253960 46998 253972
rect 48958 253960 48964 253972
rect 46992 253932 48964 253960
rect 46992 253920 46998 253932
rect 48958 253920 48964 253932
rect 49016 253920 49022 253972
rect 49050 253920 49056 253972
rect 49108 253960 49114 253972
rect 53190 253960 53196 253972
rect 49108 253932 53196 253960
rect 49108 253920 49114 253932
rect 53190 253920 53196 253932
rect 53248 253920 53254 253972
rect 144270 253920 144276 253972
rect 144328 253960 144334 253972
rect 146938 253960 146944 253972
rect 144328 253932 146944 253960
rect 144328 253920 144334 253932
rect 146938 253920 146944 253932
rect 146996 253920 147002 253972
rect 135898 252832 135904 252884
rect 135956 252872 135962 252884
rect 144270 252872 144276 252884
rect 135956 252844 144276 252872
rect 135956 252832 135962 252844
rect 144270 252832 144276 252844
rect 144328 252832 144334 252884
rect 51810 252560 51816 252612
rect 51868 252600 51874 252612
rect 53098 252600 53104 252612
rect 51868 252572 53104 252600
rect 51868 252560 51874 252572
rect 53098 252560 53104 252572
rect 53156 252560 53162 252612
rect 50338 250656 50344 250708
rect 50396 250696 50402 250708
rect 51810 250696 51816 250708
rect 50396 250668 51816 250696
rect 50396 250656 50402 250668
rect 51810 250656 51816 250668
rect 51868 250656 51874 250708
rect 45186 249772 45192 249824
rect 45244 249812 45250 249824
rect 46934 249812 46940 249824
rect 45244 249784 46940 249812
rect 45244 249772 45250 249784
rect 46934 249772 46940 249784
rect 46992 249772 46998 249824
rect 46566 245624 46572 245676
rect 46624 245664 46630 245676
rect 47578 245664 47584 245676
rect 46624 245636 47584 245664
rect 46624 245624 46630 245636
rect 47578 245624 47584 245636
rect 47636 245624 47642 245676
rect 195974 245624 195980 245676
rect 196032 245664 196038 245676
rect 197998 245664 198004 245676
rect 196032 245636 198004 245664
rect 196032 245624 196038 245636
rect 197998 245624 198004 245636
rect 198056 245624 198062 245676
rect 46934 244264 46940 244316
rect 46992 244304 46998 244316
rect 49050 244304 49056 244316
rect 46992 244276 49056 244304
rect 46992 244264 46998 244276
rect 49050 244264 49056 244276
rect 49108 244264 49114 244316
rect 413278 244264 413284 244316
rect 413336 244304 413342 244316
rect 579982 244304 579988 244316
rect 413336 244276 579988 244304
rect 413336 244264 413342 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 396534 243516 396540 243568
rect 396592 243556 396598 243568
rect 396902 243556 396908 243568
rect 396592 243528 396908 243556
rect 396592 243516 396598 243528
rect 396902 243516 396908 243528
rect 396960 243516 396966 243568
rect 133598 243040 133604 243092
rect 133656 243080 133662 243092
rect 135898 243080 135904 243092
rect 133656 243052 135904 243080
rect 133656 243040 133662 243052
rect 135898 243040 135904 243052
rect 135956 243040 135962 243092
rect 124122 242156 124128 242208
rect 124180 242196 124186 242208
rect 133598 242196 133604 242208
rect 124180 242168 133604 242196
rect 124180 242156 124186 242168
rect 133598 242156 133604 242168
rect 133656 242156 133662 242208
rect 46842 240796 46848 240848
rect 46900 240836 46906 240848
rect 124122 240836 124128 240848
rect 46900 240808 124128 240836
rect 46900 240796 46906 240808
rect 124122 240796 124128 240808
rect 124180 240796 124186 240848
rect 45646 240728 45652 240780
rect 45704 240768 45710 240780
rect 195974 240768 195980 240780
rect 45704 240740 195980 240768
rect 45704 240728 45710 240740
rect 195974 240728 195980 240740
rect 196032 240728 196038 240780
rect 45830 240524 45836 240576
rect 45888 240564 45894 240576
rect 50338 240564 50344 240576
rect 45888 240536 50344 240564
rect 45888 240524 45894 240536
rect 50338 240524 50344 240536
rect 50396 240524 50402 240576
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 5166 240224 5172 240236
rect 2832 240196 5172 240224
rect 2832 240184 2838 240196
rect 5166 240184 5172 240196
rect 5224 240184 5230 240236
rect 395338 240048 395344 240100
rect 395396 240088 395402 240100
rect 396534 240088 396540 240100
rect 395396 240060 396540 240088
rect 395396 240048 395402 240060
rect 396534 240048 396540 240060
rect 396592 240048 396598 240100
rect 45278 239844 45284 239896
rect 45336 239884 45342 239896
rect 46566 239884 46572 239896
rect 45336 239856 46572 239884
rect 45336 239844 45342 239856
rect 46566 239844 46572 239856
rect 46624 239844 46630 239896
rect 44818 239776 44824 239828
rect 44876 239816 44882 239828
rect 46842 239816 46848 239828
rect 44876 239788 46848 239816
rect 44876 239776 44882 239788
rect 46842 239776 46848 239788
rect 46900 239776 46906 239828
rect 45462 239708 45468 239760
rect 45520 239748 45526 239760
rect 46750 239748 46756 239760
rect 45520 239720 46756 239748
rect 45520 239708 45526 239720
rect 46750 239708 46756 239720
rect 46808 239708 46814 239760
rect 396534 238824 396540 238876
rect 396592 238824 396598 238876
rect 45370 238756 45376 238808
rect 45428 238796 45434 238808
rect 45646 238796 45652 238808
rect 45428 238768 45652 238796
rect 45428 238756 45434 238768
rect 45646 238756 45652 238768
rect 45704 238756 45710 238808
rect 396552 238796 396580 238824
rect 396046 238768 396580 238796
rect 396046 238728 396074 238768
rect 396534 238728 396540 238740
rect 396046 238700 396540 238728
rect 396534 238688 396540 238700
rect 396592 238688 396598 238740
rect 45738 233112 45744 233164
rect 45796 233152 45802 233164
rect 105814 233152 105820 233164
rect 45796 233124 105820 233152
rect 45796 233112 45802 233124
rect 105814 233112 105820 233124
rect 105872 233112 105878 233164
rect 44818 232976 44824 233028
rect 44876 233016 44882 233028
rect 45646 233016 45652 233028
rect 44876 232988 45652 233016
rect 44876 232976 44882 232988
rect 45646 232976 45652 232988
rect 45704 232976 45710 233028
rect 45462 232364 45468 232416
rect 45520 232404 45526 232416
rect 45738 232404 45744 232416
rect 45520 232376 45744 232404
rect 45520 232364 45526 232376
rect 45738 232364 45744 232376
rect 45796 232364 45802 232416
rect 45830 232364 45836 232416
rect 45888 232404 45894 232416
rect 48314 232404 48320 232416
rect 45888 232376 48320 232404
rect 45888 232364 45894 232376
rect 48314 232364 48320 232376
rect 48372 232364 48378 232416
rect 45370 232296 45376 232348
rect 45428 232336 45434 232348
rect 46842 232336 46848 232348
rect 45428 232308 46848 232336
rect 45428 232296 45434 232308
rect 46842 232296 46848 232308
rect 46900 232296 46906 232348
rect 394694 232092 394700 232144
rect 394752 232132 394758 232144
rect 396534 232132 396540 232144
rect 394752 232104 396540 232132
rect 394752 232092 394758 232104
rect 396534 232092 396540 232104
rect 396592 232092 396598 232144
rect 105814 231956 105820 232008
rect 105872 231996 105878 232008
rect 117958 231996 117964 232008
rect 105872 231968 117964 231996
rect 105872 231956 105878 231968
rect 117958 231956 117964 231968
rect 118016 231956 118022 232008
rect 396534 231956 396540 232008
rect 396592 231996 396598 232008
rect 396902 231996 396908 232008
rect 396592 231968 396908 231996
rect 396592 231956 396598 231968
rect 396902 231956 396908 231968
rect 396960 231956 396966 232008
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 580074 231860 580080 231872
rect 394016 231832 580080 231860
rect 394016 231820 394022 231832
rect 580074 231820 580080 231832
rect 580132 231820 580138 231872
rect 45738 231752 45744 231804
rect 45796 231792 45802 231804
rect 50614 231792 50620 231804
rect 45796 231764 50620 231792
rect 45796 231752 45802 231764
rect 50614 231752 50620 231764
rect 50672 231752 50678 231804
rect 3326 231140 3332 231192
rect 3384 231180 3390 231192
rect 179414 231180 179420 231192
rect 3384 231152 179420 231180
rect 3384 231140 3390 231152
rect 179414 231140 179420 231152
rect 179472 231140 179478 231192
rect 4062 231072 4068 231124
rect 4120 231112 4126 231124
rect 180794 231112 180800 231124
rect 4120 231084 180800 231112
rect 4120 231072 4126 231084
rect 180794 231072 180800 231084
rect 180852 231072 180858 231124
rect 45278 231004 45284 231056
rect 45336 231044 45342 231056
rect 159358 231044 159364 231056
rect 45336 231016 159364 231044
rect 45336 231004 45342 231016
rect 159358 231004 159364 231016
rect 159416 231004 159422 231056
rect 48314 230936 48320 230988
rect 48372 230976 48378 230988
rect 72418 230976 72424 230988
rect 48372 230948 72424 230976
rect 48372 230936 48378 230948
rect 72418 230936 72424 230948
rect 72476 230936 72482 230988
rect 45186 230460 45192 230512
rect 45244 230500 45250 230512
rect 46934 230500 46940 230512
rect 45244 230472 46940 230500
rect 45244 230460 45250 230472
rect 46934 230460 46940 230472
rect 46992 230460 46998 230512
rect 46842 230392 46848 230444
rect 46900 230432 46906 230444
rect 49602 230432 49608 230444
rect 46900 230404 49608 230432
rect 46900 230392 46906 230404
rect 49602 230392 49608 230404
rect 49660 230392 49666 230444
rect 45646 230324 45652 230376
rect 45704 230364 45710 230376
rect 51534 230364 51540 230376
rect 45704 230336 51540 230364
rect 45704 230324 45710 230336
rect 51534 230324 51540 230336
rect 51592 230324 51598 230376
rect 392670 229780 392676 229832
rect 392728 229820 392734 229832
rect 396626 229820 396632 229832
rect 392728 229792 396632 229820
rect 392728 229780 392734 229792
rect 396626 229780 396632 229792
rect 396684 229780 396690 229832
rect 117958 229712 117964 229764
rect 118016 229752 118022 229764
rect 131758 229752 131764 229764
rect 118016 229724 131764 229752
rect 118016 229712 118022 229724
rect 131758 229712 131764 229724
rect 131816 229712 131822 229764
rect 390922 229508 390928 229560
rect 390980 229548 390986 229560
rect 394694 229548 394700 229560
rect 390980 229520 394700 229548
rect 390980 229508 390986 229520
rect 394694 229508 394700 229520
rect 394752 229508 394758 229560
rect 157978 228420 157984 228472
rect 158036 228460 158042 228472
rect 266538 228460 266544 228472
rect 158036 228432 266544 228460
rect 158036 228420 158042 228432
rect 266538 228420 266544 228432
rect 266596 228420 266602 228472
rect 266998 228420 267004 228472
rect 267056 228460 267062 228472
rect 356514 228460 356520 228472
rect 267056 228432 356520 228460
rect 267056 228420 267062 228432
rect 356514 228420 356520 228432
rect 356572 228420 356578 228472
rect 118786 228352 118792 228404
rect 118844 228392 118850 228404
rect 580718 228392 580724 228404
rect 118844 228364 580724 228392
rect 118844 228352 118850 228364
rect 580718 228352 580724 228364
rect 580776 228352 580782 228404
rect 50614 227808 50620 227860
rect 50672 227848 50678 227860
rect 56502 227848 56508 227860
rect 50672 227820 56508 227848
rect 50672 227808 50678 227820
rect 56502 227808 56508 227820
rect 56560 227808 56566 227860
rect 2866 227740 2872 227792
rect 2924 227780 2930 227792
rect 138658 227780 138664 227792
rect 2924 227752 138664 227780
rect 2924 227740 2930 227752
rect 138658 227740 138664 227752
rect 138716 227740 138722 227792
rect 49694 227468 49700 227520
rect 49752 227508 49758 227520
rect 52362 227508 52368 227520
rect 49752 227480 52368 227508
rect 49752 227468 49758 227480
rect 52362 227468 52368 227480
rect 52420 227468 52426 227520
rect 72418 226992 72424 227044
rect 72476 227032 72482 227044
rect 77938 227032 77944 227044
rect 72476 227004 77944 227032
rect 72476 226992 72482 227004
rect 77938 226992 77944 227004
rect 77996 226992 78002 227044
rect 377306 226992 377312 227044
rect 377364 227032 377370 227044
rect 396534 227032 396540 227044
rect 377364 227004 396540 227032
rect 377364 226992 377370 227004
rect 396534 226992 396540 227004
rect 396592 226992 396598 227044
rect 384390 226856 384396 226908
rect 384448 226896 384454 226908
rect 390922 226896 390928 226908
rect 384448 226868 390928 226896
rect 384448 226856 384454 226868
rect 390922 226856 390928 226868
rect 390980 226856 390986 226908
rect 46934 225564 46940 225616
rect 46992 225604 46998 225616
rect 57882 225604 57888 225616
rect 46992 225576 57888 225604
rect 46992 225564 46998 225576
rect 57882 225564 57888 225576
rect 57940 225564 57946 225616
rect 56502 225224 56508 225276
rect 56560 225264 56566 225276
rect 57238 225264 57244 225276
rect 56560 225236 57244 225264
rect 56560 225224 56566 225236
rect 57238 225224 57244 225236
rect 57296 225224 57302 225276
rect 381538 224612 381544 224664
rect 381596 224652 381602 224664
rect 384390 224652 384396 224664
rect 381596 224624 384396 224652
rect 381596 224612 381602 224624
rect 384390 224612 384396 224624
rect 384448 224612 384454 224664
rect 51534 223592 51540 223644
rect 51592 223632 51598 223644
rect 51592 223604 55214 223632
rect 51592 223592 51598 223604
rect 55186 223564 55214 223604
rect 55858 223564 55864 223576
rect 55186 223536 55864 223564
rect 55858 223524 55864 223536
rect 55916 223524 55922 223576
rect 52454 223456 52460 223508
rect 52512 223496 52518 223508
rect 56042 223496 56048 223508
rect 52512 223468 56048 223496
rect 52512 223456 52518 223468
rect 56042 223456 56048 223468
rect 56100 223456 56106 223508
rect 57882 222844 57888 222896
rect 57940 222884 57946 222896
rect 65702 222884 65708 222896
rect 57940 222856 65708 222884
rect 57940 222844 57946 222856
rect 65702 222844 65708 222856
rect 65760 222844 65766 222896
rect 57238 222164 57244 222216
rect 57296 222204 57302 222216
rect 57296 222176 58020 222204
rect 57296 222164 57302 222176
rect 57992 222136 58020 222176
rect 60642 222136 60648 222148
rect 57992 222108 60648 222136
rect 60642 222096 60648 222108
rect 60700 222096 60706 222148
rect 44910 220804 44916 220856
rect 44968 220844 44974 220856
rect 47578 220844 47584 220856
rect 44968 220816 47584 220844
rect 44968 220804 44974 220816
rect 47578 220804 47584 220816
rect 47636 220804 47642 220856
rect 56042 220736 56048 220788
rect 56100 220776 56106 220788
rect 56962 220776 56968 220788
rect 56100 220748 56968 220776
rect 56100 220736 56106 220748
rect 56962 220736 56968 220748
rect 57020 220736 57026 220788
rect 65702 220736 65708 220788
rect 65760 220776 65766 220788
rect 69382 220776 69388 220788
rect 65760 220748 69388 220776
rect 65760 220736 65766 220748
rect 69382 220736 69388 220748
rect 69440 220736 69446 220788
rect 394050 220736 394056 220788
rect 394108 220776 394114 220788
rect 396442 220776 396448 220788
rect 394108 220748 396448 220776
rect 394108 220736 394114 220748
rect 396442 220736 396448 220748
rect 396500 220736 396506 220788
rect 368934 220056 368940 220108
rect 368992 220096 368998 220108
rect 377306 220096 377312 220108
rect 368992 220068 377312 220096
rect 368992 220056 368998 220068
rect 377306 220056 377312 220068
rect 377364 220056 377370 220108
rect 77938 218696 77944 218748
rect 77996 218736 78002 218748
rect 87506 218736 87512 218748
rect 77996 218708 87512 218736
rect 77996 218696 78002 218708
rect 87506 218696 87512 218708
rect 87564 218696 87570 218748
rect 69382 218016 69388 218068
rect 69440 218056 69446 218068
rect 69440 218028 70440 218056
rect 69440 218016 69446 218028
rect 70412 217988 70440 218028
rect 118694 218016 118700 218068
rect 118752 218056 118758 218068
rect 580074 218056 580080 218068
rect 118752 218028 580080 218056
rect 118752 218016 118758 218028
rect 580074 218016 580080 218028
rect 580132 218016 580138 218068
rect 71958 217988 71964 218000
rect 70412 217960 71964 217988
rect 71958 217948 71964 217960
rect 72016 217948 72022 218000
rect 45094 217268 45100 217320
rect 45152 217308 45158 217320
rect 53834 217308 53840 217320
rect 45152 217280 53840 217308
rect 45152 217268 45158 217280
rect 53834 217268 53840 217280
rect 53892 217268 53898 217320
rect 380158 216656 380164 216708
rect 380216 216696 380222 216708
rect 381538 216696 381544 216708
rect 380216 216668 381544 216696
rect 380216 216656 380222 216668
rect 381538 216656 381544 216668
rect 381596 216656 381602 216708
rect 45002 216588 45008 216640
rect 45060 216628 45066 216640
rect 46198 216628 46204 216640
rect 45060 216600 46204 216628
rect 45060 216588 45066 216600
rect 46198 216588 46204 216600
rect 46256 216588 46262 216640
rect 56962 216452 56968 216504
rect 57020 216492 57026 216504
rect 59630 216492 59636 216504
rect 57020 216464 59636 216492
rect 57020 216452 57026 216464
rect 59630 216452 59636 216464
rect 59688 216452 59694 216504
rect 71958 215296 71964 215348
rect 72016 215336 72022 215348
rect 72016 215308 74534 215336
rect 72016 215296 72022 215308
rect 74506 215268 74534 215308
rect 76558 215268 76564 215280
rect 74506 215240 76564 215268
rect 76558 215228 76564 215240
rect 76616 215228 76622 215280
rect 53834 214548 53840 214600
rect 53892 214588 53898 214600
rect 77938 214588 77944 214600
rect 53892 214560 77944 214588
rect 53892 214548 53898 214560
rect 77938 214548 77944 214560
rect 77996 214548 78002 214600
rect 358722 214548 358728 214600
rect 358780 214588 358786 214600
rect 368934 214588 368940 214600
rect 358780 214560 368940 214588
rect 358780 214548 358786 214560
rect 368934 214548 368940 214560
rect 368992 214548 368998 214600
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 179506 213976 179512 213988
rect 3384 213948 179512 213976
rect 3384 213936 3390 213948
rect 179506 213936 179512 213948
rect 179564 213936 179570 213988
rect 60734 213868 60740 213920
rect 60792 213908 60798 213920
rect 63494 213908 63500 213920
rect 60792 213880 63500 213908
rect 60792 213868 60798 213880
rect 63494 213868 63500 213880
rect 63552 213868 63558 213920
rect 59630 213188 59636 213240
rect 59688 213228 59694 213240
rect 68278 213228 68284 213240
rect 59688 213200 68284 213228
rect 59688 213188 59694 213200
rect 68278 213188 68284 213200
rect 68336 213188 68342 213240
rect 47578 212440 47584 212492
rect 47636 212480 47642 212492
rect 52454 212480 52460 212492
rect 47636 212452 52460 212480
rect 47636 212440 47642 212452
rect 52454 212440 52460 212452
rect 52512 212440 52518 212492
rect 55858 212440 55864 212492
rect 55916 212480 55922 212492
rect 59262 212480 59268 212492
rect 55916 212452 59268 212480
rect 55916 212440 55922 212452
rect 59262 212440 59268 212452
rect 59320 212440 59326 212492
rect 344094 211760 344100 211812
rect 344152 211800 344158 211812
rect 358722 211800 358728 211812
rect 344152 211772 358728 211800
rect 344152 211760 344158 211772
rect 358722 211760 358728 211772
rect 358780 211760 358786 211812
rect 63494 211012 63500 211064
rect 63552 211052 63558 211064
rect 65886 211052 65892 211064
rect 63552 211024 65892 211052
rect 63552 211012 63558 211024
rect 65886 211012 65892 211024
rect 65944 211012 65950 211064
rect 87506 209788 87512 209840
rect 87564 209828 87570 209840
rect 95878 209828 95884 209840
rect 87564 209800 95884 209828
rect 87564 209788 87570 209800
rect 95878 209788 95884 209800
rect 95936 209788 95942 209840
rect 159358 209788 159364 209840
rect 159416 209828 159422 209840
rect 162118 209828 162124 209840
rect 159416 209800 162124 209828
rect 159416 209788 159422 209800
rect 162118 209788 162124 209800
rect 162176 209788 162182 209840
rect 392578 209788 392584 209840
rect 392636 209828 392642 209840
rect 394050 209828 394056 209840
rect 392636 209800 394056 209828
rect 392636 209788 392642 209800
rect 394050 209788 394056 209800
rect 394108 209788 394114 209840
rect 59262 209108 59268 209160
rect 59320 209148 59326 209160
rect 62114 209148 62120 209160
rect 59320 209120 62120 209148
rect 59320 209108 59326 209120
rect 62114 209108 62120 209120
rect 62172 209108 62178 209160
rect 46198 208972 46204 209024
rect 46256 209012 46262 209024
rect 48774 209012 48780 209024
rect 46256 208984 48780 209012
rect 46256 208972 46262 208984
rect 48774 208972 48780 208984
rect 48832 208972 48838 209024
rect 68278 208904 68284 208956
rect 68336 208944 68342 208956
rect 75546 208944 75552 208956
rect 68336 208916 75552 208944
rect 68336 208904 68342 208916
rect 75546 208904 75552 208916
rect 75604 208904 75610 208956
rect 52454 208632 52460 208684
rect 52512 208672 52518 208684
rect 55858 208672 55864 208684
rect 52512 208644 55864 208672
rect 52512 208632 52518 208644
rect 55858 208632 55864 208644
rect 55916 208632 55922 208684
rect 65886 208360 65892 208412
rect 65944 208400 65950 208412
rect 65944 208372 67680 208400
rect 65944 208360 65950 208372
rect 67652 208332 67680 208372
rect 376754 208360 376760 208412
rect 376812 208400 376818 208412
rect 380158 208400 380164 208412
rect 376812 208372 380164 208400
rect 376812 208360 376818 208372
rect 380158 208360 380164 208372
rect 380216 208360 380222 208412
rect 71682 208332 71688 208344
rect 67652 208304 71688 208332
rect 71682 208292 71688 208304
rect 71740 208292 71746 208344
rect 341518 207000 341524 207052
rect 341576 207040 341582 207052
rect 344094 207040 344100 207052
rect 341576 207012 344100 207040
rect 341576 207000 341582 207012
rect 344094 207000 344100 207012
rect 344152 207000 344158 207052
rect 389174 207000 389180 207052
rect 389232 207040 389238 207052
rect 392670 207040 392676 207052
rect 389232 207012 392676 207040
rect 389232 207000 389238 207012
rect 392670 207000 392676 207012
rect 392728 207000 392734 207052
rect 62114 205640 62120 205692
rect 62172 205680 62178 205692
rect 62172 205652 64874 205680
rect 62172 205640 62178 205652
rect 48774 205572 48780 205624
rect 48832 205612 48838 205624
rect 56410 205612 56416 205624
rect 48832 205584 56416 205612
rect 48832 205572 48838 205584
rect 56410 205572 56416 205584
rect 56468 205572 56474 205624
rect 64846 205612 64874 205652
rect 189718 205640 189724 205692
rect 189776 205680 189782 205692
rect 580074 205680 580080 205692
rect 189776 205652 580080 205680
rect 189776 205640 189782 205652
rect 580074 205640 580080 205652
rect 580132 205640 580138 205692
rect 66438 205612 66444 205624
rect 64846 205584 66444 205612
rect 66438 205572 66444 205584
rect 66496 205572 66502 205624
rect 76558 205368 76564 205420
rect 76616 205408 76622 205420
rect 78306 205408 78312 205420
rect 76616 205380 78312 205408
rect 76616 205368 76622 205380
rect 78306 205368 78312 205380
rect 78364 205368 78370 205420
rect 377674 204892 377680 204944
rect 377732 204932 377738 204944
rect 389174 204932 389180 204944
rect 377732 204904 389180 204932
rect 377732 204892 377738 204904
rect 389174 204892 389180 204904
rect 389232 204892 389238 204944
rect 71774 204212 71780 204264
rect 71832 204252 71838 204264
rect 73798 204252 73804 204264
rect 71832 204224 73804 204252
rect 71832 204212 71838 204224
rect 73798 204212 73804 204224
rect 73856 204212 73862 204264
rect 56410 202920 56416 202972
rect 56468 202960 56474 202972
rect 62114 202960 62120 202972
rect 56468 202932 62120 202960
rect 56468 202920 56474 202932
rect 62114 202920 62120 202932
rect 62172 202920 62178 202972
rect 373994 202240 374000 202292
rect 374052 202280 374058 202292
rect 377674 202280 377680 202292
rect 374052 202252 377680 202280
rect 374052 202240 374058 202252
rect 377674 202240 377680 202252
rect 377732 202240 377738 202292
rect 147766 202104 147772 202156
rect 147824 202144 147830 202156
rect 176654 202144 176660 202156
rect 147824 202116 176660 202144
rect 147824 202104 147830 202116
rect 176654 202104 176660 202116
rect 176712 202104 176718 202156
rect 3326 201832 3332 201884
rect 3384 201872 3390 201884
rect 7558 201872 7564 201884
rect 3384 201844 7564 201872
rect 3384 201832 3390 201844
rect 7558 201832 7564 201844
rect 7616 201832 7622 201884
rect 62114 201424 62120 201476
rect 62172 201464 62178 201476
rect 64230 201464 64236 201476
rect 62172 201436 64236 201464
rect 62172 201424 62178 201436
rect 64230 201424 64236 201436
rect 64288 201424 64294 201476
rect 66438 201424 66444 201476
rect 66496 201464 66502 201476
rect 69658 201464 69664 201476
rect 66496 201436 69664 201464
rect 66496 201424 66502 201436
rect 69658 201424 69664 201436
rect 69716 201424 69722 201476
rect 75546 201424 75552 201476
rect 75604 201464 75610 201476
rect 76558 201464 76564 201476
rect 75604 201436 76564 201464
rect 75604 201424 75610 201436
rect 76558 201424 76564 201436
rect 76616 201424 76622 201476
rect 77938 201424 77944 201476
rect 77996 201464 78002 201476
rect 80698 201464 80704 201476
rect 77996 201436 80704 201464
rect 77996 201424 78002 201436
rect 80698 201424 80704 201436
rect 80756 201424 80762 201476
rect 78306 201356 78312 201408
rect 78364 201396 78370 201408
rect 79962 201396 79968 201408
rect 78364 201368 79968 201396
rect 78364 201356 78370 201368
rect 79962 201356 79968 201368
rect 80020 201356 80026 201408
rect 375374 201288 375380 201340
rect 375432 201328 375438 201340
rect 376754 201328 376760 201340
rect 375432 201300 376760 201328
rect 375432 201288 375438 201300
rect 376754 201288 376760 201300
rect 376812 201288 376818 201340
rect 155954 199384 155960 199436
rect 156012 199424 156018 199436
rect 296714 199424 296720 199436
rect 156012 199396 296720 199424
rect 156012 199384 156018 199396
rect 296714 199384 296720 199396
rect 296772 199384 296778 199436
rect 351178 199384 351184 199436
rect 351236 199424 351242 199436
rect 373994 199424 374000 199436
rect 351236 199396 374000 199424
rect 351236 199384 351242 199396
rect 373994 199384 374000 199396
rect 374052 199384 374058 199436
rect 338758 198704 338764 198756
rect 338816 198744 338822 198756
rect 341518 198744 341524 198756
rect 338816 198716 341524 198744
rect 338816 198704 338822 198716
rect 341518 198704 341524 198716
rect 341576 198704 341582 198756
rect 73798 198228 73804 198280
rect 73856 198268 73862 198280
rect 75546 198268 75552 198280
rect 73856 198240 75552 198268
rect 73856 198228 73862 198240
rect 75546 198228 75552 198240
rect 75604 198228 75610 198280
rect 148962 197956 148968 198008
rect 149020 197996 149026 198008
rect 207014 197996 207020 198008
rect 149020 197968 207020 197996
rect 149020 197956 149026 197968
rect 207014 197956 207020 197968
rect 207072 197956 207078 198008
rect 154482 197412 154488 197464
rect 154540 197452 154546 197464
rect 155954 197452 155960 197464
rect 154540 197424 155960 197452
rect 154540 197412 154546 197424
rect 155954 197412 155960 197424
rect 156012 197412 156018 197464
rect 79962 197344 79968 197396
rect 80020 197384 80026 197396
rect 80020 197356 81480 197384
rect 80020 197344 80026 197356
rect 81452 197316 81480 197356
rect 84838 197316 84844 197328
rect 81452 197288 84844 197316
rect 84838 197276 84844 197288
rect 84896 197276 84902 197328
rect 152734 197276 152740 197328
rect 152792 197316 152798 197328
rect 157978 197316 157984 197328
rect 152792 197288 157984 197316
rect 152792 197276 152798 197288
rect 157978 197276 157984 197288
rect 158036 197276 158042 197328
rect 138658 196732 138664 196784
rect 138716 196772 138722 196784
rect 164234 196772 164240 196784
rect 138716 196744 164240 196772
rect 138716 196732 138722 196744
rect 164234 196732 164240 196744
rect 164292 196732 164298 196784
rect 151170 196664 151176 196716
rect 151228 196704 151234 196716
rect 235994 196704 236000 196716
rect 151228 196676 236000 196704
rect 151228 196664 151234 196676
rect 235994 196664 236000 196676
rect 236052 196664 236058 196716
rect 155954 196596 155960 196648
rect 156012 196636 156018 196648
rect 327074 196636 327080 196648
rect 156012 196608 327080 196636
rect 156012 196596 156018 196608
rect 327074 196596 327080 196608
rect 327132 196596 327138 196648
rect 162118 196460 162124 196512
rect 162176 196500 162182 196512
rect 164142 196500 164148 196512
rect 162176 196472 164148 196500
rect 162176 196460 162182 196472
rect 164142 196460 164148 196472
rect 164200 196460 164206 196512
rect 367094 196460 367100 196512
rect 367152 196500 367158 196512
rect 375374 196500 375380 196512
rect 367152 196472 375380 196500
rect 367152 196460 367158 196472
rect 375374 196460 375380 196472
rect 375432 196460 375438 196512
rect 56594 195916 56600 195968
rect 56652 195956 56658 195968
rect 138106 195956 138112 195968
rect 56652 195928 138112 195956
rect 56652 195916 56658 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 160094 195916 160100 195968
rect 160152 195956 160158 195968
rect 386414 195956 386420 195968
rect 160152 195928 386420 195956
rect 160152 195916 160158 195928
rect 386414 195916 386420 195928
rect 386472 195916 386478 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 157610 195848 157616 195900
rect 157668 195888 157674 195900
rect 266998 195888 267004 195900
rect 157668 195860 267004 195888
rect 157668 195848 157674 195860
rect 266998 195848 267004 195860
rect 267056 195848 267062 195900
rect 75546 194624 75552 194676
rect 75604 194664 75610 194676
rect 76650 194664 76656 194676
rect 75604 194636 76656 194664
rect 75604 194624 75610 194636
rect 76650 194624 76656 194636
rect 76708 194624 76714 194676
rect 115934 194556 115940 194608
rect 115992 194596 115998 194608
rect 140774 194596 140780 194608
rect 115992 194568 140780 194596
rect 115992 194556 115998 194568
rect 140774 194556 140780 194568
rect 140832 194556 140838 194608
rect 164142 194488 164148 194540
rect 164200 194528 164206 194540
rect 167638 194528 167644 194540
rect 164200 194500 167644 194528
rect 164200 194488 164206 194500
rect 167638 194488 167644 194500
rect 167696 194488 167702 194540
rect 504450 191836 504456 191888
rect 504508 191876 504514 191888
rect 579798 191876 579804 191888
rect 504508 191848 579804 191876
rect 504508 191836 504514 191848
rect 579798 191836 579804 191848
rect 579856 191836 579862 191888
rect 55858 191768 55864 191820
rect 55916 191808 55922 191820
rect 64138 191808 64144 191820
rect 55916 191780 64144 191808
rect 55916 191768 55922 191780
rect 64138 191768 64144 191780
rect 64196 191768 64202 191820
rect 144454 190476 144460 190528
rect 144512 190516 144518 190528
rect 144512 190488 145052 190516
rect 144512 190476 144518 190488
rect 145024 190324 145052 190488
rect 362218 190476 362224 190528
rect 362276 190516 362282 190528
rect 367002 190516 367008 190528
rect 362276 190488 367008 190516
rect 362276 190476 362282 190488
rect 367002 190476 367008 190488
rect 367060 190476 367066 190528
rect 145006 190272 145012 190324
rect 145064 190272 145070 190324
rect 64230 189728 64236 189780
rect 64288 189768 64294 189780
rect 69750 189768 69756 189780
rect 64288 189740 69756 189768
rect 64288 189728 64294 189740
rect 69750 189728 69756 189740
rect 69808 189728 69814 189780
rect 144638 189048 144644 189100
rect 144696 189088 144702 189100
rect 145006 189088 145012 189100
rect 144696 189060 145012 189088
rect 144696 189048 144702 189060
rect 145006 189048 145012 189060
rect 145064 189048 145070 189100
rect 76558 188164 76564 188216
rect 76616 188204 76622 188216
rect 78582 188204 78588 188216
rect 76616 188176 78588 188204
rect 76616 188164 76622 188176
rect 78582 188164 78588 188176
rect 78640 188164 78646 188216
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 115198 187728 115204 187740
rect 3384 187700 115204 187728
rect 3384 187688 3390 187700
rect 115198 187688 115204 187700
rect 115256 187688 115262 187740
rect 335998 187688 336004 187740
rect 336056 187728 336062 187740
rect 338758 187728 338764 187740
rect 336056 187700 338764 187728
rect 336056 187688 336062 187700
rect 338758 187688 338764 187700
rect 338816 187688 338822 187740
rect 76650 187348 76656 187400
rect 76708 187388 76714 187400
rect 79962 187388 79968 187400
rect 76708 187360 79968 187388
rect 76708 187348 76714 187360
rect 79962 187348 79968 187360
rect 80020 187348 80026 187400
rect 84838 186940 84844 186992
rect 84896 186980 84902 186992
rect 86218 186980 86224 186992
rect 84896 186952 86224 186980
rect 84896 186940 84902 186952
rect 86218 186940 86224 186952
rect 86276 186940 86282 186992
rect 69658 185988 69664 186040
rect 69716 186028 69722 186040
rect 71038 186028 71044 186040
rect 69716 186000 71044 186028
rect 69716 185988 69722 186000
rect 71038 185988 71044 186000
rect 71096 185988 71102 186040
rect 159542 185852 159548 185904
rect 159600 185852 159606 185904
rect 159560 185552 159588 185852
rect 159910 185552 159916 185564
rect 159560 185524 159916 185552
rect 159910 185512 159916 185524
rect 159968 185512 159974 185564
rect 79962 184832 79968 184884
rect 80020 184872 80026 184884
rect 81434 184872 81440 184884
rect 80020 184844 81440 184872
rect 80020 184832 80026 184844
rect 81434 184832 81440 184844
rect 81492 184832 81498 184884
rect 78674 184764 78680 184816
rect 78732 184804 78738 184816
rect 80790 184804 80796 184816
rect 78732 184776 80796 184804
rect 78732 184764 78738 184776
rect 80790 184764 80796 184776
rect 80848 184764 80854 184816
rect 390554 183472 390560 183524
rect 390612 183512 390618 183524
rect 392578 183512 392584 183524
rect 390612 183484 392584 183512
rect 390612 183472 390618 183484
rect 392578 183472 392584 183484
rect 392636 183472 392642 183524
rect 131758 183404 131764 183456
rect 131816 183444 131822 183456
rect 133966 183444 133972 183456
rect 131816 183416 133972 183444
rect 131816 183404 131822 183416
rect 133966 183404 133972 183416
rect 134024 183404 134030 183456
rect 81434 182180 81440 182232
rect 81492 182220 81498 182232
rect 81492 182192 84194 182220
rect 81492 182180 81498 182192
rect 84166 182152 84194 182192
rect 86310 182152 86316 182164
rect 84166 182124 86316 182152
rect 86310 182112 86316 182124
rect 86368 182112 86374 182164
rect 144638 181092 144644 181144
rect 144696 181092 144702 181144
rect 144656 181064 144684 181092
rect 151906 181064 151912 181076
rect 144656 181036 151912 181064
rect 151906 181024 151912 181036
rect 151964 181024 151970 181076
rect 159910 180684 159916 180736
rect 159968 180684 159974 180736
rect 140056 180288 140774 180316
rect 121454 180140 121460 180192
rect 121512 180180 121518 180192
rect 136358 180180 136364 180192
rect 121512 180152 136364 180180
rect 121512 180140 121518 180152
rect 136358 180140 136364 180152
rect 136416 180140 136422 180192
rect 133966 180072 133972 180124
rect 134024 180112 134030 180124
rect 140056 180112 140084 180288
rect 134024 180084 140084 180112
rect 134024 180072 134030 180084
rect 140746 179432 140774 180288
rect 159928 180124 159956 180684
rect 159910 180072 159916 180124
rect 159968 180072 159974 180124
rect 151906 179460 151912 179512
rect 151964 179500 151970 179512
rect 153930 179500 153936 179512
rect 151964 179472 153936 179500
rect 151964 179460 151970 179472
rect 153930 179460 153936 179472
rect 153988 179460 153994 179512
rect 149054 179432 149060 179444
rect 140746 179404 149060 179432
rect 149054 179392 149060 179404
rect 149112 179392 149118 179444
rect 154390 179392 154396 179444
rect 154448 179432 154454 179444
rect 157794 179432 157800 179444
rect 154448 179404 157800 179432
rect 154448 179392 154454 179404
rect 157794 179392 157800 179404
rect 157852 179392 157858 179444
rect 158622 179392 158628 179444
rect 158680 179432 158686 179444
rect 169754 179432 169760 179444
rect 158680 179404 169760 179432
rect 158680 179392 158686 179404
rect 169754 179392 169760 179404
rect 169812 179392 169818 179444
rect 136726 178780 136732 178832
rect 136784 178780 136790 178832
rect 122834 178644 122840 178696
rect 122892 178684 122898 178696
rect 136450 178684 136456 178696
rect 122892 178656 136456 178684
rect 122892 178644 122898 178656
rect 136450 178644 136456 178656
rect 136508 178644 136514 178696
rect 136358 178372 136364 178424
rect 136416 178412 136422 178424
rect 136744 178412 136772 178780
rect 136416 178384 136772 178412
rect 136416 178372 136422 178384
rect 71038 178304 71044 178356
rect 71096 178344 71102 178356
rect 72418 178344 72424 178356
rect 71096 178316 72424 178344
rect 71096 178304 71102 178316
rect 72418 178304 72424 178316
rect 72476 178304 72482 178356
rect 330018 177964 330024 178016
rect 330076 178004 330082 178016
rect 335998 178004 336004 178016
rect 330076 177976 336004 178004
rect 330076 177964 330082 177976
rect 335998 177964 336004 177976
rect 336056 177964 336062 178016
rect 134978 177760 134984 177812
rect 135036 177800 135042 177812
rect 136634 177800 136640 177812
rect 135036 177772 136640 177800
rect 135036 177760 135042 177772
rect 136634 177760 136640 177772
rect 136692 177760 136698 177812
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 136450 177324 136456 177336
rect 124272 177296 136456 177324
rect 124272 177284 124278 177296
rect 136450 177284 136456 177296
rect 136508 177284 136514 177336
rect 135254 177216 135260 177268
rect 135312 177256 135318 177268
rect 136542 177256 136548 177268
rect 135312 177228 136548 177256
rect 135312 177216 135318 177228
rect 136542 177216 136548 177228
rect 136600 177216 136606 177268
rect 159910 176400 159916 176452
rect 159968 176400 159974 176452
rect 126974 176128 126980 176180
rect 127032 176168 127038 176180
rect 134978 176168 134984 176180
rect 127032 176140 134984 176168
rect 127032 176128 127038 176140
rect 134978 176128 134984 176140
rect 135036 176128 135042 176180
rect 125594 175992 125600 176044
rect 125652 176032 125658 176044
rect 136358 176032 136364 176044
rect 125652 176004 136364 176032
rect 125652 175992 125658 176004
rect 136358 175992 136364 176004
rect 136416 175992 136422 176044
rect 144086 175992 144092 176044
rect 144144 176032 144150 176044
rect 149330 176032 149336 176044
rect 144144 176004 149336 176032
rect 144144 175992 144150 176004
rect 149330 175992 149336 176004
rect 149388 175992 149394 176044
rect 159928 176032 159956 176400
rect 159192 176004 159956 176032
rect 69750 175924 69756 175976
rect 69808 175964 69814 175976
rect 92474 175964 92480 175976
rect 69808 175936 92480 175964
rect 69808 175924 69814 175936
rect 92474 175924 92480 175936
rect 92532 175924 92538 175976
rect 118878 175924 118884 175976
rect 118936 175964 118942 175976
rect 118936 175936 142154 175964
rect 118936 175924 118942 175936
rect 142126 175760 142154 175936
rect 158686 175936 159036 175964
rect 144454 175788 144460 175840
rect 144512 175828 144518 175840
rect 149974 175828 149980 175840
rect 144512 175800 149980 175828
rect 144512 175788 144518 175800
rect 149974 175788 149980 175800
rect 150032 175788 150038 175840
rect 154408 175800 157334 175828
rect 142126 175732 144914 175760
rect 144886 175420 144914 175732
rect 154408 175432 154436 175800
rect 157306 175692 157334 175800
rect 158162 175720 158168 175772
rect 158220 175760 158226 175772
rect 158686 175760 158714 175936
rect 158220 175732 158714 175760
rect 159008 175760 159036 175936
rect 159192 175908 159220 176004
rect 165062 175924 165068 175976
rect 165120 175964 165126 175976
rect 580074 175964 580080 175976
rect 165120 175936 580080 175964
rect 165120 175924 165126 175936
rect 580074 175924 580080 175936
rect 580132 175924 580138 175976
rect 159174 175856 159180 175908
rect 159232 175856 159238 175908
rect 165154 175856 165160 175908
rect 165212 175896 165218 175908
rect 166994 175896 167000 175908
rect 165212 175868 167000 175896
rect 165212 175856 165218 175868
rect 166994 175856 167000 175868
rect 167052 175856 167058 175908
rect 163498 175760 163504 175772
rect 159008 175732 163504 175760
rect 158220 175720 158226 175732
rect 163498 175720 163504 175732
rect 163556 175720 163562 175772
rect 163590 175692 163596 175704
rect 157306 175664 163596 175692
rect 163590 175652 163596 175664
rect 163648 175652 163654 175704
rect 153930 175420 153936 175432
rect 144886 175392 153936 175420
rect 153930 175380 153936 175392
rect 153988 175380 153994 175432
rect 154390 175380 154396 175432
rect 154448 175380 154454 175432
rect 159174 175420 159180 175432
rect 157306 175392 159180 175420
rect 155494 175244 155500 175296
rect 155552 175284 155558 175296
rect 157306 175284 157334 175392
rect 159174 175380 159180 175392
rect 159232 175380 159238 175432
rect 155552 175256 157334 175284
rect 155552 175244 155558 175256
rect 128354 175176 128360 175228
rect 128412 175216 128418 175228
rect 135254 175216 135260 175228
rect 128412 175188 135260 175216
rect 128412 175176 128418 175188
rect 135254 175176 135260 175188
rect 135312 175176 135318 175228
rect 385678 175176 385684 175228
rect 385736 175216 385742 175228
rect 390462 175216 390468 175228
rect 385736 175188 390468 175216
rect 385736 175176 385742 175188
rect 390462 175176 390468 175188
rect 390520 175176 390526 175228
rect 141602 174768 141608 174820
rect 141660 174808 141666 174820
rect 146478 174808 146484 174820
rect 141660 174780 146484 174808
rect 141660 174768 141666 174780
rect 146478 174768 146484 174780
rect 146536 174768 146542 174820
rect 149054 174768 149060 174820
rect 149112 174808 149118 174820
rect 149112 174780 153194 174808
rect 149112 174768 149118 174780
rect 143074 174700 143080 174752
rect 143132 174740 143138 174752
rect 143132 174712 144914 174740
rect 143132 174700 143138 174712
rect 144886 174604 144914 174712
rect 152366 174700 152372 174752
rect 152424 174700 152430 174752
rect 153166 174740 153194 174780
rect 162486 174740 162492 174752
rect 153166 174712 162492 174740
rect 162486 174700 162492 174712
rect 162544 174700 162550 174752
rect 152384 174672 152412 174700
rect 156506 174672 156512 174684
rect 152384 174644 156512 174672
rect 156506 174632 156512 174644
rect 156564 174632 156570 174684
rect 161474 174604 161480 174616
rect 144886 174576 161480 174604
rect 161474 174564 161480 174576
rect 161532 174564 161538 174616
rect 155494 174536 155500 174548
rect 141712 174508 155500 174536
rect 135898 174360 135904 174412
rect 135956 174400 135962 174412
rect 141712 174400 141740 174508
rect 155494 174496 155500 174508
rect 155552 174496 155558 174548
rect 135956 174372 141740 174400
rect 135956 174360 135962 174372
rect 146478 174292 146484 174344
rect 146536 174332 146542 174344
rect 146536 174304 165476 174332
rect 146536 174292 146542 174304
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 137370 173924 137376 173936
rect 133932 173896 137376 173924
rect 133932 173884 133938 173896
rect 137370 173884 137376 173896
rect 137428 173884 137434 173936
rect 86310 173816 86316 173868
rect 86368 173856 86374 173868
rect 87966 173856 87972 173868
rect 86368 173828 87972 173856
rect 86368 173816 86374 173828
rect 87966 173816 87972 173828
rect 88024 173816 88030 173868
rect 165448 172984 165476 174304
rect 327718 174088 327724 174140
rect 327776 174128 327782 174140
rect 330018 174128 330024 174140
rect 327776 174100 330024 174128
rect 327776 174088 327782 174100
rect 330018 174088 330024 174100
rect 330076 174088 330082 174140
rect 167638 173816 167644 173868
rect 167696 173856 167702 173868
rect 169110 173856 169116 173868
rect 167696 173828 169116 173856
rect 167696 173816 167702 173828
rect 169110 173816 169116 173828
rect 169168 173816 169174 173868
rect 149330 172932 149336 172984
rect 149388 172972 149394 172984
rect 150434 172972 150440 172984
rect 149388 172944 150440 172972
rect 149388 172932 149394 172944
rect 150434 172932 150440 172944
rect 150492 172932 150498 172984
rect 165430 172932 165436 172984
rect 165488 172932 165494 172984
rect 131114 172524 131120 172576
rect 131172 172564 131178 172576
rect 136542 172564 136548 172576
rect 131172 172536 136548 172564
rect 131172 172524 131178 172536
rect 136542 172524 136548 172536
rect 136600 172524 136606 172576
rect 359826 172456 359832 172508
rect 359884 172496 359890 172508
rect 362218 172496 362224 172508
rect 359884 172468 362224 172496
rect 359884 172456 359890 172468
rect 362218 172456 362224 172468
rect 362276 172456 362282 172508
rect 138014 172116 138020 172168
rect 138072 172156 138078 172168
rect 140774 172156 140780 172168
rect 138072 172128 140780 172156
rect 138072 172116 138078 172128
rect 140774 172116 140780 172128
rect 140832 172116 140838 172168
rect 64138 171776 64144 171828
rect 64196 171816 64202 171828
rect 69934 171816 69940 171828
rect 64196 171788 69940 171816
rect 64196 171776 64202 171788
rect 69934 171776 69940 171788
rect 69992 171776 69998 171828
rect 135254 171640 135260 171692
rect 135312 171680 135318 171692
rect 138658 171680 138664 171692
rect 135312 171652 138664 171680
rect 135312 171640 135318 171652
rect 138658 171640 138664 171652
rect 138716 171640 138722 171692
rect 92474 171368 92480 171420
rect 92532 171408 92538 171420
rect 94498 171408 94504 171420
rect 92532 171380 94504 171408
rect 92532 171368 92538 171380
rect 94498 171368 94504 171380
rect 94556 171368 94562 171420
rect 132494 171096 132500 171148
rect 132552 171136 132558 171148
rect 136726 171136 136732 171148
rect 132552 171108 136732 171136
rect 132552 171096 132558 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 162854 169940 162860 169992
rect 162912 169980 162918 169992
rect 163498 169980 163504 169992
rect 162912 169952 163504 169980
rect 162912 169940 162918 169952
rect 163498 169940 163504 169952
rect 163556 169940 163562 169992
rect 87966 169804 87972 169856
rect 88024 169844 88030 169856
rect 88978 169844 88984 169856
rect 88024 169816 88984 169844
rect 88024 169804 88030 169816
rect 88978 169804 88984 169816
rect 89036 169804 89042 169856
rect 169110 169736 169116 169788
rect 169168 169776 169174 169788
rect 170398 169776 170404 169788
rect 169168 169748 170404 169776
rect 169168 169736 169174 169748
rect 170398 169736 170404 169748
rect 170456 169736 170462 169788
rect 346302 169736 346308 169788
rect 346360 169776 346366 169788
rect 351178 169776 351184 169788
rect 346360 169748 351184 169776
rect 346360 169736 346366 169748
rect 351178 169736 351184 169748
rect 351236 169736 351242 169788
rect 86218 168852 86224 168904
rect 86276 168892 86282 168904
rect 88334 168892 88340 168904
rect 86276 168864 88340 168892
rect 86276 168852 86282 168864
rect 88334 168852 88340 168864
rect 88392 168852 88398 168904
rect 69934 168240 69940 168292
rect 69992 168280 69998 168292
rect 77202 168280 77208 168292
rect 69992 168252 77208 168280
rect 69992 168240 69998 168252
rect 77202 168240 77208 168252
rect 77260 168240 77266 168292
rect 80698 168240 80704 168292
rect 80756 168280 80762 168292
rect 86862 168280 86868 168292
rect 80756 168252 86868 168280
rect 80756 168240 80762 168252
rect 86862 168240 86868 168252
rect 86920 168240 86926 168292
rect 80790 167016 80796 167068
rect 80848 167056 80854 167068
rect 82078 167056 82084 167068
rect 80848 167028 82084 167056
rect 80848 167016 80854 167028
rect 82078 167016 82084 167028
rect 82136 167016 82142 167068
rect 163590 166336 163596 166388
rect 163648 166336 163654 166388
rect 163608 166184 163636 166336
rect 163590 166132 163596 166184
rect 163648 166132 163654 166184
rect 340138 166064 340144 166116
rect 340196 166104 340202 166116
rect 346302 166104 346308 166116
rect 340196 166076 346308 166104
rect 340196 166064 340202 166076
rect 346302 166064 346308 166076
rect 346360 166064 346366 166116
rect 188338 165588 188344 165640
rect 188396 165628 188402 165640
rect 580074 165628 580080 165640
rect 188396 165600 580080 165628
rect 188396 165588 188402 165600
rect 580074 165588 580080 165600
rect 580132 165588 580138 165640
rect 88334 165520 88340 165572
rect 88392 165560 88398 165572
rect 90358 165560 90364 165572
rect 88392 165532 90364 165560
rect 88392 165520 88398 165532
rect 90358 165520 90364 165532
rect 90416 165520 90422 165572
rect 356698 165316 356704 165368
rect 356756 165356 356762 165368
rect 359826 165356 359832 165368
rect 356756 165328 359832 165356
rect 356756 165316 356762 165328
rect 359826 165316 359832 165328
rect 359884 165316 359890 165368
rect 77202 164840 77208 164892
rect 77260 164880 77266 164892
rect 85206 164880 85212 164892
rect 77260 164852 85212 164880
rect 77260 164840 77266 164852
rect 85206 164840 85212 164852
rect 85264 164840 85270 164892
rect 118970 164840 118976 164892
rect 119028 164880 119034 164892
rect 580810 164880 580816 164892
rect 119028 164852 580816 164880
rect 119028 164840 119034 164852
rect 580810 164840 580816 164852
rect 580868 164840 580874 164892
rect 86862 164160 86868 164212
rect 86920 164200 86926 164212
rect 91554 164200 91560 164212
rect 86920 164172 91560 164200
rect 86920 164160 86926 164172
rect 91554 164160 91560 164172
rect 91612 164160 91618 164212
rect 155218 164160 155224 164212
rect 155276 164200 155282 164212
rect 160094 164200 160100 164212
rect 155276 164172 160100 164200
rect 155276 164160 155282 164172
rect 160094 164160 160100 164172
rect 160152 164160 160158 164212
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 181254 162908 181260 162920
rect 3384 162880 181260 162908
rect 3384 162868 3390 162880
rect 181254 162868 181260 162880
rect 181312 162868 181318 162920
rect 85206 162800 85212 162852
rect 85264 162840 85270 162852
rect 91738 162840 91744 162852
rect 85264 162812 91744 162840
rect 85264 162800 85270 162812
rect 91738 162800 91744 162812
rect 91796 162800 91802 162852
rect 20070 162120 20076 162172
rect 20128 162160 20134 162172
rect 182910 162160 182916 162172
rect 20128 162132 182916 162160
rect 20128 162120 20134 162132
rect 182910 162120 182916 162132
rect 182968 162120 182974 162172
rect 324314 161440 324320 161492
rect 324372 161480 324378 161492
rect 327718 161480 327724 161492
rect 324372 161452 327724 161480
rect 324372 161440 324378 161452
rect 327718 161440 327724 161452
rect 327776 161440 327782 161492
rect 170398 160692 170404 160744
rect 170456 160732 170462 160744
rect 173894 160732 173900 160744
rect 170456 160704 173900 160732
rect 170456 160692 170462 160704
rect 173894 160692 173900 160704
rect 173952 160692 173958 160744
rect 72418 160420 72424 160472
rect 72476 160460 72482 160472
rect 76742 160460 76748 160472
rect 72476 160432 76748 160460
rect 72476 160420 72482 160432
rect 76742 160420 76748 160432
rect 76800 160420 76806 160472
rect 94498 160080 94504 160132
rect 94556 160120 94562 160132
rect 94556 160092 96660 160120
rect 94556 160080 94562 160092
rect 96632 160052 96660 160092
rect 163682 160080 163688 160132
rect 163740 160120 163746 160132
rect 166258 160120 166264 160132
rect 163740 160092 166264 160120
rect 163740 160080 163746 160092
rect 166258 160080 166264 160092
rect 166316 160080 166322 160132
rect 382274 160080 382280 160132
rect 382332 160120 382338 160132
rect 385678 160120 385684 160132
rect 382332 160092 385684 160120
rect 382332 160080 382338 160092
rect 385678 160080 385684 160092
rect 385736 160080 385742 160132
rect 98638 160052 98644 160064
rect 96632 160024 98644 160052
rect 98638 160012 98644 160024
rect 98696 160012 98702 160064
rect 91554 159332 91560 159384
rect 91612 159372 91618 159384
rect 98178 159372 98184 159384
rect 91612 159344 98184 159372
rect 91612 159332 91618 159344
rect 98178 159332 98184 159344
rect 98236 159332 98242 159384
rect 319898 158720 319904 158772
rect 319956 158760 319962 158772
rect 324314 158760 324320 158772
rect 319956 158732 324320 158760
rect 319956 158720 319962 158732
rect 324314 158720 324320 158732
rect 324372 158720 324378 158772
rect 82078 158040 82084 158092
rect 82136 158080 82142 158092
rect 83458 158080 83464 158092
rect 82136 158052 83464 158080
rect 82136 158040 82142 158052
rect 83458 158040 83464 158052
rect 83516 158040 83522 158092
rect 160094 158040 160100 158092
rect 160152 158080 160158 158092
rect 166350 158080 166356 158092
rect 160152 158052 166356 158080
rect 160152 158040 160158 158052
rect 166350 158040 166356 158052
rect 166408 158040 166414 158092
rect 119062 157972 119068 158024
rect 119120 158012 119126 158024
rect 580166 158012 580172 158024
rect 119120 157984 580172 158012
rect 119120 157972 119126 157984
rect 580166 157972 580172 157984
rect 580224 157972 580230 158024
rect 173894 157632 173900 157684
rect 173952 157672 173958 157684
rect 175918 157672 175924 157684
rect 173952 157644 175924 157672
rect 173952 157632 173958 157644
rect 175918 157632 175924 157644
rect 175976 157632 175982 157684
rect 356698 155972 356704 155984
rect 354646 155944 356704 155972
rect 76742 155864 76748 155916
rect 76800 155904 76806 155916
rect 79318 155904 79324 155916
rect 76800 155876 79324 155904
rect 76800 155864 76806 155876
rect 79318 155864 79324 155876
rect 79376 155864 79382 155916
rect 353938 155864 353944 155916
rect 353996 155904 354002 155916
rect 354646 155904 354674 155944
rect 356698 155932 356704 155944
rect 356756 155932 356762 155984
rect 382182 155972 382188 155984
rect 376772 155944 382188 155972
rect 353996 155876 354674 155904
rect 353996 155864 354002 155876
rect 374638 155864 374644 155916
rect 374696 155904 374702 155916
rect 376772 155904 376800 155944
rect 382182 155932 382188 155944
rect 382240 155932 382246 155984
rect 374696 155876 376800 155904
rect 374696 155864 374702 155876
rect 303982 155184 303988 155236
rect 304040 155224 304046 155236
rect 319898 155224 319904 155236
rect 304040 155196 319904 155224
rect 304040 155184 304046 155196
rect 319898 155184 319904 155196
rect 319956 155184 319962 155236
rect 322198 155184 322204 155236
rect 322256 155224 322262 155236
rect 340138 155224 340144 155236
rect 322256 155196 340144 155224
rect 322256 155184 322262 155196
rect 340138 155184 340144 155196
rect 340196 155184 340202 155236
rect 98178 153144 98184 153196
rect 98236 153184 98242 153196
rect 102778 153184 102784 153196
rect 98236 153156 102784 153184
rect 98236 153144 98242 153156
rect 102778 153144 102784 153156
rect 102836 153144 102842 153196
rect 301498 152804 301504 152856
rect 301556 152844 301562 152856
rect 303982 152844 303988 152856
rect 301556 152816 303988 152844
rect 301556 152804 301562 152816
rect 303982 152804 303988 152816
rect 304040 152804 304046 152856
rect 180058 151784 180064 151836
rect 180116 151824 180122 151836
rect 579982 151824 579988 151836
rect 180116 151796 579988 151824
rect 180116 151784 180122 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 88978 150424 88984 150476
rect 89036 150464 89042 150476
rect 89036 150436 91140 150464
rect 89036 150424 89042 150436
rect 91112 150396 91140 150436
rect 372614 150424 372620 150476
rect 372672 150464 372678 150476
rect 374638 150464 374644 150476
rect 372672 150436 374644 150464
rect 372672 150424 372678 150436
rect 374638 150424 374644 150436
rect 374696 150424 374702 150476
rect 94774 150396 94780 150408
rect 91112 150368 94780 150396
rect 94774 150356 94780 150368
rect 94832 150356 94838 150408
rect 3234 149676 3240 149728
rect 3292 149716 3298 149728
rect 22922 149716 22928 149728
rect 3292 149688 22928 149716
rect 3292 149676 3298 149688
rect 22922 149676 22928 149688
rect 22980 149676 22986 149728
rect 91738 148316 91744 148368
rect 91796 148356 91802 148368
rect 109678 148356 109684 148368
rect 91796 148328 109684 148356
rect 91796 148316 91802 148328
rect 109678 148316 109684 148328
rect 109736 148316 109742 148368
rect 134058 147636 134064 147688
rect 134116 147676 134122 147688
rect 135898 147676 135904 147688
rect 134116 147648 135904 147676
rect 134116 147636 134122 147648
rect 135898 147636 135904 147648
rect 135956 147636 135962 147688
rect 45554 146956 45560 147008
rect 45612 146996 45618 147008
rect 48958 146996 48964 147008
rect 45612 146968 48964 146996
rect 45612 146956 45618 146968
rect 48958 146956 48964 146968
rect 49016 146956 49022 147008
rect 166350 146956 166356 147008
rect 166408 146996 166414 147008
rect 168374 146996 168380 147008
rect 166408 146968 168380 146996
rect 166408 146956 166414 146968
rect 168374 146956 168380 146968
rect 168432 146956 168438 147008
rect 166258 146888 166264 146940
rect 166316 146928 166322 146940
rect 180150 146928 180156 146940
rect 166316 146900 180156 146928
rect 166316 146888 166322 146900
rect 180150 146888 180156 146900
rect 180208 146888 180214 146940
rect 94774 146276 94780 146328
rect 94832 146316 94838 146328
rect 94832 146288 95280 146316
rect 94832 146276 94838 146288
rect 95252 146248 95280 146288
rect 371878 146276 371884 146328
rect 371936 146316 371942 146328
rect 372614 146316 372620 146328
rect 371936 146288 372620 146316
rect 371936 146276 371942 146288
rect 372614 146276 372620 146288
rect 372672 146276 372678 146328
rect 97258 146248 97264 146260
rect 95252 146220 97264 146248
rect 97258 146208 97264 146220
rect 97316 146208 97322 146260
rect 141694 146208 141700 146260
rect 141752 146248 141758 146260
rect 142430 146248 142436 146260
rect 141752 146220 142436 146248
rect 141752 146208 141758 146220
rect 142430 146208 142436 146220
rect 142488 146208 142494 146260
rect 350534 144780 350540 144832
rect 350592 144820 350598 144832
rect 353938 144820 353944 144832
rect 350592 144792 353944 144820
rect 350592 144780 350598 144792
rect 353938 144780 353944 144792
rect 353996 144780 354002 144832
rect 33778 144440 33784 144492
rect 33836 144480 33842 144492
rect 182634 144480 182640 144492
rect 33836 144452 182640 144480
rect 33836 144440 33842 144452
rect 182634 144440 182640 144452
rect 182692 144440 182698 144492
rect 10410 144372 10416 144424
rect 10468 144412 10474 144424
rect 182542 144412 182548 144424
rect 10468 144384 182548 144412
rect 10468 144372 10474 144384
rect 182542 144372 182548 144384
rect 182600 144372 182606 144424
rect 6178 144304 6184 144356
rect 6236 144344 6242 144356
rect 182266 144344 182272 144356
rect 6236 144316 182272 144344
rect 6236 144304 6242 144316
rect 182266 144304 182272 144316
rect 182324 144304 182330 144356
rect 118326 144236 118332 144288
rect 118384 144276 118390 144288
rect 398190 144276 398196 144288
rect 118384 144248 398196 144276
rect 118384 144236 118390 144248
rect 398190 144236 398196 144248
rect 398248 144236 398254 144288
rect 118234 144168 118240 144220
rect 118292 144208 118298 144220
rect 398098 144208 398104 144220
rect 118292 144180 398104 144208
rect 118292 144168 118298 144180
rect 398098 144168 398104 144180
rect 398156 144168 398162 144220
rect 98638 143488 98644 143540
rect 98696 143528 98702 143540
rect 100938 143528 100944 143540
rect 98696 143500 100944 143528
rect 98696 143488 98702 143500
rect 100938 143488 100944 143500
rect 100996 143488 101002 143540
rect 146478 143488 146484 143540
rect 146536 143528 146542 143540
rect 148042 143528 148048 143540
rect 146536 143500 148048 143528
rect 146536 143488 146542 143500
rect 148042 143488 148048 143500
rect 148100 143488 148106 143540
rect 153470 143488 153476 143540
rect 153528 143528 153534 143540
rect 158990 143528 158996 143540
rect 153528 143500 158996 143528
rect 153528 143488 153534 143500
rect 158990 143488 158996 143500
rect 159048 143488 159054 143540
rect 147674 143420 147680 143472
rect 147732 143460 147738 143472
rect 149606 143460 149612 143472
rect 147732 143432 149612 143460
rect 147732 143420 147738 143432
rect 149606 143420 149612 143432
rect 149664 143420 149670 143472
rect 152458 143420 152464 143472
rect 152516 143460 152522 143472
rect 157426 143460 157432 143472
rect 152516 143432 157432 143460
rect 152516 143420 152522 143432
rect 157426 143420 157432 143432
rect 157484 143420 157490 143472
rect 137738 143352 137744 143404
rect 137796 143392 137802 143404
rect 139578 143392 139584 143404
rect 137796 143364 139584 143392
rect 137796 143352 137802 143364
rect 139578 143352 139584 143364
rect 139636 143352 139642 143404
rect 163590 143148 163596 143200
rect 163648 143188 163654 143200
rect 174630 143188 174636 143200
rect 163648 143160 174636 143188
rect 163648 143148 163654 143160
rect 174630 143148 174636 143160
rect 174688 143148 174694 143200
rect 150526 143080 150532 143132
rect 150584 143120 150590 143132
rect 154574 143120 154580 143132
rect 150584 143092 154580 143120
rect 150584 143080 150590 143092
rect 154574 143080 154580 143092
rect 154632 143080 154638 143132
rect 164510 143080 164516 143132
rect 164568 143120 164574 143132
rect 176194 143120 176200 143132
rect 164568 143092 176200 143120
rect 164568 143080 164574 143092
rect 176194 143080 176200 143092
rect 176252 143080 176258 143132
rect 122834 143012 122840 143064
rect 122892 143052 122898 143064
rect 134058 143052 134064 143064
rect 122892 143024 134064 143052
rect 122892 143012 122898 143024
rect 134058 143012 134064 143024
rect 134116 143012 134122 143064
rect 144454 143012 144460 143064
rect 144512 143052 144518 143064
rect 160554 143052 160560 143064
rect 144512 143024 160560 143052
rect 144512 143012 144518 143024
rect 160554 143012 160560 143024
rect 160612 143012 160618 143064
rect 163498 143012 163504 143064
rect 163556 143052 163562 143064
rect 178034 143052 178040 143064
rect 163556 143024 178040 143052
rect 163556 143012 163562 143024
rect 178034 143012 178040 143024
rect 178092 143012 178098 143064
rect 118510 142944 118516 142996
rect 118568 142984 118574 142996
rect 398374 142984 398380 142996
rect 118568 142956 398380 142984
rect 118568 142944 118574 142956
rect 398374 142944 398380 142956
rect 398432 142944 398438 142996
rect 118418 142876 118424 142928
rect 118476 142916 118482 142928
rect 398282 142916 398288 142928
rect 118476 142888 398288 142916
rect 118476 142876 118482 142888
rect 398282 142876 398288 142888
rect 398340 142876 398346 142928
rect 102778 142808 102784 142860
rect 102836 142848 102842 142860
rect 108298 142848 108304 142860
rect 102836 142820 108304 142848
rect 102836 142808 102842 142820
rect 108298 142808 108304 142820
rect 108356 142808 108362 142860
rect 120718 142808 120724 142860
rect 120776 142848 120782 142860
rect 477494 142848 477500 142860
rect 120776 142820 477500 142848
rect 120776 142808 120782 142820
rect 477494 142808 477500 142820
rect 477552 142808 477558 142860
rect 140682 142128 140688 142180
rect 140740 142168 140746 142180
rect 142154 142168 142160 142180
rect 140740 142140 142160 142168
rect 140740 142128 140746 142140
rect 142154 142128 142160 142140
rect 142212 142128 142218 142180
rect 149514 142128 149520 142180
rect 149572 142168 149578 142180
rect 152734 142168 152740 142180
rect 149572 142140 152740 142168
rect 149572 142128 149578 142140
rect 152734 142128 152740 142140
rect 152792 142128 152798 142180
rect 157334 142128 157340 142180
rect 157392 142168 157398 142180
rect 163682 142168 163688 142180
rect 157392 142140 163688 142168
rect 157392 142128 157398 142140
rect 163682 142128 163688 142140
rect 163740 142128 163746 142180
rect 175918 142128 175924 142180
rect 175976 142168 175982 142180
rect 175976 142140 176700 142168
rect 175976 142128 175982 142140
rect 176672 142100 176700 142140
rect 181162 142100 181168 142112
rect 176672 142072 181168 142100
rect 181162 142060 181168 142072
rect 181220 142060 181226 142112
rect 40034 141652 40040 141704
rect 40092 141692 40098 141704
rect 180978 141692 180984 141704
rect 40092 141664 180984 141692
rect 40092 141652 40098 141664
rect 180978 141652 180984 141664
rect 181036 141652 181042 141704
rect 4890 141584 4896 141636
rect 4948 141624 4954 141636
rect 182450 141624 182456 141636
rect 4948 141596 182456 141624
rect 4948 141584 4954 141596
rect 182450 141584 182456 141596
rect 182508 141584 182514 141636
rect 118142 141516 118148 141568
rect 118200 141556 118206 141568
rect 542354 141556 542360 141568
rect 118200 141528 542360 141556
rect 118200 141516 118206 141528
rect 542354 141516 542360 141528
rect 542412 141516 542418 141568
rect 119246 141448 119252 141500
rect 119304 141488 119310 141500
rect 580258 141488 580264 141500
rect 119304 141460 580264 141488
rect 119304 141448 119310 141460
rect 580258 141448 580264 141460
rect 580316 141448 580322 141500
rect 119154 141380 119160 141432
rect 119212 141420 119218 141432
rect 580534 141420 580540 141432
rect 119212 141392 580540 141420
rect 119212 141380 119218 141392
rect 580534 141380 580540 141392
rect 580592 141380 580598 141432
rect 121270 140428 121276 140480
rect 121328 140468 121334 140480
rect 122834 140468 122840 140480
rect 121328 140440 122840 140468
rect 121328 140428 121334 140440
rect 122834 140428 122840 140440
rect 122892 140428 122898 140480
rect 79318 140292 79324 140344
rect 79376 140332 79382 140344
rect 82722 140332 82728 140344
rect 79376 140304 82728 140332
rect 79376 140292 79382 140304
rect 82722 140292 82728 140304
rect 82780 140292 82786 140344
rect 100938 140292 100944 140344
rect 100996 140332 101002 140344
rect 181070 140332 181076 140344
rect 100996 140304 181076 140332
rect 100996 140292 101002 140304
rect 181070 140292 181076 140304
rect 181128 140292 181134 140344
rect 10318 140224 10324 140276
rect 10376 140264 10382 140276
rect 182726 140264 182732 140276
rect 10376 140236 182732 140264
rect 10376 140224 10382 140236
rect 182726 140224 182732 140236
rect 182784 140224 182790 140276
rect 4798 140156 4804 140208
rect 4856 140196 4862 140208
rect 182358 140196 182364 140208
rect 4856 140168 182364 140196
rect 4856 140156 4862 140168
rect 182358 140156 182364 140168
rect 182416 140156 182422 140208
rect 83458 140088 83464 140140
rect 83516 140128 83522 140140
rect 85022 140128 85028 140140
rect 83516 140100 85028 140128
rect 83516 140088 83522 140100
rect 85022 140088 85028 140100
rect 85080 140088 85086 140140
rect 119982 140088 119988 140140
rect 120040 140128 120046 140140
rect 301498 140128 301504 140140
rect 120040 140100 301504 140128
rect 120040 140088 120046 140100
rect 301498 140088 301504 140100
rect 301556 140088 301562 140140
rect 118050 140020 118056 140072
rect 118108 140060 118114 140072
rect 412634 140060 412640 140072
rect 118108 140032 412640 140060
rect 118108 140020 118114 140032
rect 412634 140020 412640 140032
rect 412692 140020 412698 140072
rect 90358 139816 90364 139868
rect 90416 139856 90422 139868
rect 91462 139856 91468 139868
rect 90416 139828 91468 139856
rect 90416 139816 90422 139828
rect 91462 139816 91468 139828
rect 91520 139816 91526 139868
rect 118602 139476 118608 139528
rect 118660 139516 118666 139528
rect 178218 139516 178224 139528
rect 118660 139488 178224 139516
rect 118660 139476 118666 139488
rect 178218 139476 178224 139488
rect 178276 139476 178282 139528
rect 43438 139408 43444 139460
rect 43496 139448 43502 139460
rect 182174 139448 182180 139460
rect 43496 139420 182180 139448
rect 43496 139408 43502 139420
rect 182174 139408 182180 139420
rect 182232 139408 182238 139460
rect 369762 139408 369768 139460
rect 369820 139448 369826 139460
rect 371878 139448 371884 139460
rect 369820 139420 371884 139448
rect 369820 139408 369826 139420
rect 371878 139408 371884 139420
rect 371936 139408 371942 139460
rect 178218 139340 178224 139392
rect 178276 139380 178282 139392
rect 580166 139380 580172 139392
rect 178276 139352 580172 139380
rect 178276 139340 178282 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 4062 138660 4068 138712
rect 4120 138700 4126 138712
rect 25498 138700 25504 138712
rect 4120 138672 25504 138700
rect 4120 138660 4126 138672
rect 25498 138660 25504 138672
rect 25556 138660 25562 138712
rect 85022 138048 85028 138100
rect 85080 138088 85086 138100
rect 86218 138088 86224 138100
rect 85080 138060 86224 138088
rect 85080 138048 85086 138060
rect 86218 138048 86224 138060
rect 86276 138048 86282 138100
rect 367738 137980 367744 138032
rect 367796 138020 367802 138032
rect 369762 138020 369768 138032
rect 367796 137992 369768 138020
rect 367796 137980 367802 137992
rect 369762 137980 369768 137992
rect 369820 137980 369826 138032
rect 4062 136688 4068 136740
rect 4120 136728 4126 136740
rect 117314 136728 117320 136740
rect 4120 136700 117320 136728
rect 4120 136688 4126 136700
rect 117314 136688 117320 136700
rect 117372 136688 117378 136740
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 119338 136660 119344 136672
rect 3384 136632 119344 136660
rect 3384 136620 3390 136632
rect 119338 136620 119344 136632
rect 119396 136620 119402 136672
rect 350534 136660 350540 136672
rect 347792 136632 350540 136660
rect 345658 136552 345664 136604
rect 345716 136592 345722 136604
rect 347792 136592 347820 136632
rect 350534 136620 350540 136632
rect 350592 136620 350598 136672
rect 345716 136564 347820 136592
rect 345716 136552 345722 136564
rect 117958 136144 117964 136196
rect 118016 136184 118022 136196
rect 119982 136184 119988 136196
rect 118016 136156 119988 136184
rect 118016 136144 118022 136156
rect 119982 136144 119988 136156
rect 120040 136144 120046 136196
rect 3326 135260 3332 135312
rect 3384 135300 3390 135312
rect 117314 135300 117320 135312
rect 3384 135272 117320 135300
rect 3384 135260 3390 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 91462 135192 91468 135244
rect 91520 135232 91526 135244
rect 93762 135232 93768 135244
rect 91520 135204 93768 135232
rect 91520 135192 91526 135204
rect 93762 135192 93768 135204
rect 93820 135192 93826 135244
rect 82814 134852 82820 134904
rect 82872 134892 82878 134904
rect 85206 134892 85212 134904
rect 82872 134864 85212 134892
rect 82872 134852 82878 134864
rect 85206 134852 85212 134864
rect 85264 134852 85270 134904
rect 295978 134512 295984 134564
rect 296036 134552 296042 134564
rect 322198 134552 322204 134564
rect 296036 134524 322204 134552
rect 296036 134512 296042 134524
rect 322198 134512 322204 134524
rect 322256 134512 322262 134564
rect 3234 133900 3240 133952
rect 3292 133940 3298 133952
rect 117314 133940 117320 133952
rect 3292 133912 117320 133940
rect 3292 133900 3298 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 108298 133152 108304 133204
rect 108356 133192 108362 133204
rect 117774 133192 117780 133204
rect 108356 133164 117780 133192
rect 108356 133152 108362 133164
rect 117774 133152 117780 133164
rect 117832 133152 117838 133204
rect 25498 132404 25504 132456
rect 25556 132444 25562 132456
rect 117314 132444 117320 132456
rect 25556 132416 117320 132444
rect 25556 132404 25562 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 86218 131112 86224 131164
rect 86276 131152 86282 131164
rect 89530 131152 89536 131164
rect 86276 131124 89536 131152
rect 86276 131112 86282 131124
rect 89530 131112 89536 131124
rect 89588 131112 89594 131164
rect 180150 131112 180156 131164
rect 180208 131152 180214 131164
rect 182174 131152 182180 131164
rect 180208 131124 182180 131152
rect 180208 131112 180214 131124
rect 182174 131112 182180 131124
rect 182232 131112 182238 131164
rect 365714 131112 365720 131164
rect 365772 131152 365778 131164
rect 367738 131152 367744 131164
rect 365772 131124 367744 131152
rect 365772 131112 365778 131124
rect 367738 131112 367744 131124
rect 367796 131112 367802 131164
rect 7558 131044 7564 131096
rect 7616 131084 7622 131096
rect 117314 131084 117320 131096
rect 7616 131056 117320 131084
rect 7616 131044 7622 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 93854 130092 93860 130144
rect 93912 130132 93918 130144
rect 95602 130132 95608 130144
rect 93912 130104 95608 130132
rect 93912 130092 93918 130104
rect 95602 130092 95608 130104
rect 95660 130092 95666 130144
rect 22830 129684 22836 129736
rect 22888 129724 22894 129736
rect 117314 129724 117320 129736
rect 22888 129696 117320 129724
rect 22888 129684 22894 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 89530 129616 89536 129668
rect 89588 129656 89594 129668
rect 92382 129656 92388 129668
rect 89588 129628 92388 129656
rect 89588 129616 89594 129628
rect 92382 129616 92388 129628
rect 92440 129616 92446 129668
rect 97258 128596 97264 128648
rect 97316 128636 97322 128648
rect 99742 128636 99748 128648
rect 97316 128608 99748 128636
rect 97316 128596 97322 128608
rect 99742 128596 99748 128608
rect 99800 128596 99806 128648
rect 109678 128324 109684 128376
rect 109736 128364 109742 128376
rect 112438 128364 112444 128376
rect 109736 128336 112444 128364
rect 109736 128324 109742 128336
rect 112438 128324 112444 128336
rect 112496 128324 112502 128376
rect 22922 128256 22928 128308
rect 22980 128296 22986 128308
rect 117314 128296 117320 128308
rect 22980 128268 117320 128296
rect 22980 128256 22986 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 363598 127712 363604 127764
rect 363656 127752 363662 127764
rect 365714 127752 365720 127764
rect 363656 127724 365720 127752
rect 363656 127712 363662 127724
rect 365714 127712 365720 127724
rect 365772 127712 365778 127764
rect 22738 126896 22744 126948
rect 22796 126936 22802 126948
rect 117314 126936 117320 126948
rect 22796 126908 117320 126936
rect 22796 126896 22802 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 85206 126828 85212 126880
rect 85264 126868 85270 126880
rect 88794 126868 88800 126880
rect 85264 126840 88800 126868
rect 85264 126828 85270 126840
rect 88794 126828 88800 126840
rect 88852 126828 88858 126880
rect 182818 125604 182824 125656
rect 182876 125644 182882 125656
rect 580166 125644 580172 125656
rect 182876 125616 580172 125644
rect 182876 125604 182882 125616
rect 580166 125604 580172 125616
rect 580224 125604 580230 125656
rect 8938 125536 8944 125588
rect 8996 125576 9002 125588
rect 117314 125576 117320 125588
rect 8996 125548 117320 125576
rect 8996 125536 9002 125548
rect 117314 125536 117320 125548
rect 117372 125536 117378 125588
rect 95602 125468 95608 125520
rect 95660 125508 95666 125520
rect 97166 125508 97172 125520
rect 95660 125480 97172 125508
rect 95660 125468 95666 125480
rect 97166 125468 97172 125480
rect 97224 125468 97230 125520
rect 345658 124216 345664 124228
rect 344986 124188 345664 124216
rect 4982 124108 4988 124160
rect 5040 124148 5046 124160
rect 117314 124148 117320 124160
rect 5040 124120 117320 124148
rect 5040 124108 5046 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 342254 124108 342260 124160
rect 342312 124148 342318 124160
rect 344986 124148 345014 124188
rect 345658 124176 345664 124188
rect 345716 124176 345722 124228
rect 342312 124120 345014 124148
rect 342312 124108 342318 124120
rect 88794 124040 88800 124092
rect 88852 124080 88858 124092
rect 92382 124080 92388 124092
rect 88852 124052 92388 124080
rect 88852 124040 88858 124052
rect 92382 124040 92388 124052
rect 92440 124040 92446 124092
rect 99742 124040 99748 124092
rect 99800 124080 99806 124092
rect 102042 124080 102048 124092
rect 99800 124052 102048 124080
rect 99800 124040 99806 124052
rect 102042 124040 102048 124052
rect 102100 124040 102106 124092
rect 92474 123428 92480 123480
rect 92532 123468 92538 123480
rect 100754 123468 100760 123480
rect 92532 123440 100760 123468
rect 92532 123428 92538 123440
rect 100754 123428 100760 123440
rect 100812 123428 100818 123480
rect 24118 122748 24124 122800
rect 24176 122788 24182 122800
rect 117314 122788 117320 122800
rect 24176 122760 117320 122788
rect 24176 122748 24182 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 100754 121796 100760 121848
rect 100812 121836 100818 121848
rect 102134 121836 102140 121848
rect 100812 121808 102140 121836
rect 100812 121796 100818 121808
rect 102134 121796 102140 121808
rect 102192 121796 102198 121848
rect 92382 121728 92388 121780
rect 92440 121768 92446 121780
rect 94406 121768 94412 121780
rect 92440 121740 94412 121768
rect 92440 121728 92446 121740
rect 94406 121728 94412 121740
rect 94464 121728 94470 121780
rect 37918 121388 37924 121440
rect 37976 121428 37982 121440
rect 117314 121428 117320 121440
rect 37976 121400 117320 121428
rect 37976 121388 37982 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 97166 120844 97172 120896
rect 97224 120884 97230 120896
rect 105722 120884 105728 120896
rect 97224 120856 105728 120884
rect 97224 120844 97230 120856
rect 105722 120844 105728 120856
rect 105780 120844 105786 120896
rect 19978 120028 19984 120080
rect 20036 120068 20042 120080
rect 117314 120068 117320 120080
rect 20036 120040 117320 120068
rect 20036 120028 20042 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 102042 119960 102048 120012
rect 102100 120000 102106 120012
rect 104342 120000 104348 120012
rect 102100 119972 104348 120000
rect 102100 119960 102106 119972
rect 104342 119960 104348 119972
rect 104400 119960 104406 120012
rect 15838 118600 15844 118652
rect 15896 118640 15902 118652
rect 117314 118640 117320 118652
rect 15896 118612 117320 118640
rect 15896 118600 15902 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 117958 118600 117964 118652
rect 118016 118600 118022 118652
rect 102134 118532 102140 118584
rect 102192 118572 102198 118584
rect 104710 118572 104716 118584
rect 102192 118544 104716 118572
rect 102192 118532 102198 118544
rect 104710 118532 104716 118544
rect 104768 118532 104774 118584
rect 112438 118532 112444 118584
rect 112496 118572 112502 118584
rect 115474 118572 115480 118584
rect 112496 118544 115480 118572
rect 112496 118532 112502 118544
rect 115474 118532 115480 118544
rect 115532 118532 115538 118584
rect 104342 118396 104348 118448
rect 104400 118436 104406 118448
rect 108298 118436 108304 118448
rect 104400 118408 108304 118436
rect 104400 118396 104406 118408
rect 108298 118396 108304 118408
rect 108356 118396 108362 118448
rect 117976 118436 118004 118600
rect 118050 118436 118056 118448
rect 117976 118408 118056 118436
rect 118050 118396 118056 118408
rect 118108 118396 118114 118448
rect 94406 118260 94412 118312
rect 94464 118300 94470 118312
rect 97166 118300 97172 118312
rect 94464 118272 97172 118300
rect 94464 118260 94470 118272
rect 97166 118260 97172 118272
rect 97224 118260 97230 118312
rect 48958 117920 48964 117972
rect 49016 117960 49022 117972
rect 63494 117960 63500 117972
rect 49016 117932 63500 117960
rect 49016 117920 49022 117932
rect 63494 117920 63500 117932
rect 63552 117920 63558 117972
rect 360194 117648 360200 117700
rect 360252 117688 360258 117700
rect 363598 117688 363604 117700
rect 360252 117660 363604 117688
rect 360252 117648 360258 117660
rect 363598 117648 363604 117660
rect 363656 117648 363662 117700
rect 23474 117240 23480 117292
rect 23532 117280 23538 117292
rect 117314 117280 117320 117292
rect 23532 117252 117320 117280
rect 23532 117240 23538 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 293218 116968 293224 117020
rect 293276 117008 293282 117020
rect 295978 117008 295984 117020
rect 293276 116980 295984 117008
rect 293276 116968 293282 116980
rect 295978 116968 295984 116980
rect 296036 116968 296042 117020
rect 97166 115948 97172 116000
rect 97224 115988 97230 116000
rect 342254 115988 342260 116000
rect 97224 115960 98776 115988
rect 97224 115948 97230 115960
rect 95878 115880 95884 115932
rect 95936 115920 95942 115932
rect 98638 115920 98644 115932
rect 95936 115892 98644 115920
rect 95936 115880 95942 115892
rect 98638 115880 98644 115892
rect 98696 115880 98702 115932
rect 98748 115920 98776 115960
rect 340892 115960 342260 115988
rect 100662 115920 100668 115932
rect 98748 115892 100668 115920
rect 100662 115880 100668 115892
rect 100720 115880 100726 115932
rect 105722 115880 105728 115932
rect 105780 115920 105786 115932
rect 110322 115920 110328 115932
rect 105780 115892 110328 115920
rect 105780 115880 105786 115892
rect 110322 115880 110328 115892
rect 110380 115880 110386 115932
rect 115474 115880 115480 115932
rect 115532 115920 115538 115932
rect 117774 115920 117780 115932
rect 115532 115892 117780 115920
rect 115532 115880 115538 115892
rect 117774 115880 117780 115892
rect 117832 115880 117838 115932
rect 338758 115880 338764 115932
rect 338816 115920 338822 115932
rect 340892 115920 340920 115960
rect 342254 115948 342260 115960
rect 342312 115948 342318 116000
rect 338816 115892 340920 115920
rect 338816 115880 338822 115892
rect 358262 115064 358268 115116
rect 358320 115104 358326 115116
rect 360194 115104 360200 115116
rect 358320 115076 360200 115104
rect 358320 115064 358326 115076
rect 360194 115064 360200 115076
rect 360252 115064 360258 115116
rect 63494 114452 63500 114504
rect 63552 114492 63558 114504
rect 117314 114492 117320 114504
rect 63552 114464 117320 114492
rect 63552 114452 63558 114464
rect 117314 114452 117320 114464
rect 117372 114452 117378 114504
rect 117682 114452 117688 114504
rect 117740 114492 117746 114504
rect 120902 114492 120908 114504
rect 117740 114464 120908 114492
rect 117740 114452 117746 114464
rect 120902 114452 120908 114464
rect 120960 114452 120966 114504
rect 104710 114384 104716 114436
rect 104768 114424 104774 114436
rect 107930 114424 107936 114436
rect 104768 114396 107936 114424
rect 104768 114384 104774 114396
rect 107930 114384 107936 114396
rect 107988 114384 107994 114436
rect 351914 113772 351920 113824
rect 351972 113812 351978 113824
rect 358262 113812 358268 113824
rect 351972 113784 358268 113812
rect 351972 113772 351978 113784
rect 358262 113772 358268 113784
rect 358320 113772 358326 113824
rect 110322 113092 110328 113144
rect 110380 113132 110386 113144
rect 117314 113132 117320 113144
rect 110380 113104 117320 113132
rect 110380 113092 110386 113104
rect 117314 113092 117320 113104
rect 117372 113092 117378 113144
rect 336734 111868 336740 111920
rect 336792 111908 336798 111920
rect 338758 111908 338764 111920
rect 336792 111880 338764 111908
rect 336792 111868 336798 111880
rect 338758 111868 338764 111880
rect 338816 111868 338822 111920
rect 349154 111868 349160 111920
rect 349212 111908 349218 111920
rect 351914 111908 351920 111920
rect 349212 111880 351920 111908
rect 349212 111868 349218 111880
rect 351914 111868 351920 111880
rect 351972 111868 351978 111920
rect 180150 111800 180156 111852
rect 180208 111840 180214 111852
rect 580166 111840 580172 111852
rect 180208 111812 580172 111840
rect 180208 111800 180214 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 43438 111772 43444 111784
rect 3200 111744 43444 111772
rect 3200 111732 3206 111744
rect 43438 111732 43444 111744
rect 43496 111732 43502 111784
rect 100662 111732 100668 111784
rect 100720 111772 100726 111784
rect 117314 111772 117320 111784
rect 100720 111744 117320 111772
rect 100720 111732 100726 111744
rect 117314 111732 117320 111744
rect 117372 111732 117378 111784
rect 183278 111732 183284 111784
rect 183336 111772 183342 111784
rect 336734 111772 336740 111784
rect 183336 111744 336740 111772
rect 183336 111732 183342 111744
rect 336734 111732 336740 111744
rect 336792 111732 336798 111784
rect 107930 110440 107936 110492
rect 107988 110480 107994 110492
rect 349154 110480 349160 110492
rect 107988 110452 113174 110480
rect 107988 110440 107994 110452
rect 113146 110412 113174 110452
rect 348436 110452 349160 110480
rect 117314 110412 117320 110424
rect 113146 110384 117320 110412
rect 117314 110372 117320 110384
rect 117372 110372 117378 110424
rect 183462 110372 183468 110424
rect 183520 110412 183526 110424
rect 348436 110412 348464 110452
rect 349154 110440 349160 110452
rect 349212 110440 349218 110492
rect 183520 110384 348464 110412
rect 183520 110372 183526 110384
rect 183370 108944 183376 108996
rect 183428 108984 183434 108996
rect 410518 108984 410524 108996
rect 183428 108956 410524 108984
rect 183428 108944 183434 108956
rect 410518 108944 410524 108956
rect 410576 108944 410582 108996
rect 183462 106224 183468 106276
rect 183520 106264 183526 106276
rect 409138 106264 409144 106276
rect 183520 106236 409144 106264
rect 183520 106224 183526 106236
rect 409138 106224 409144 106236
rect 409196 106224 409202 106276
rect 183462 104796 183468 104848
rect 183520 104836 183526 104848
rect 407758 104836 407764 104848
rect 183520 104808 407764 104836
rect 183520 104796 183526 104808
rect 407758 104796 407764 104808
rect 407816 104796 407822 104848
rect 183462 103436 183468 103488
rect 183520 103476 183526 103488
rect 406378 103476 406384 103488
rect 183520 103448 406384 103476
rect 183520 103436 183526 103448
rect 406378 103436 406384 103448
rect 406436 103436 406442 103488
rect 183462 102076 183468 102128
rect 183520 102116 183526 102128
rect 404998 102116 405004 102128
rect 183520 102088 405004 102116
rect 183520 102076 183526 102088
rect 404998 102076 405004 102088
rect 405056 102076 405062 102128
rect 98638 100648 98644 100700
rect 98696 100688 98702 100700
rect 100754 100688 100760 100700
rect 98696 100660 100760 100688
rect 98696 100648 98702 100660
rect 100754 100648 100760 100660
rect 100812 100648 100818 100700
rect 183462 100648 183468 100700
rect 183520 100688 183526 100700
rect 403618 100688 403624 100700
rect 183520 100660 403624 100688
rect 183520 100648 183526 100660
rect 403618 100648 403624 100660
rect 403676 100648 403682 100700
rect 183462 99288 183468 99340
rect 183520 99328 183526 99340
rect 400858 99328 400864 99340
rect 183520 99300 400864 99328
rect 183520 99288 183526 99300
rect 400858 99288 400864 99300
rect 400916 99288 400922 99340
rect 108298 98676 108304 98728
rect 108356 98716 108362 98728
rect 109678 98716 109684 98728
rect 108356 98688 109684 98716
rect 108356 98676 108362 98688
rect 109678 98676 109684 98688
rect 109736 98676 109742 98728
rect 117774 97928 117780 97980
rect 117832 97968 117838 97980
rect 120902 97968 120908 97980
rect 117832 97940 120908 97968
rect 117832 97928 117838 97940
rect 120902 97928 120908 97940
rect 120960 97928 120966 97980
rect 183462 97928 183468 97980
rect 183520 97968 183526 97980
rect 399478 97968 399484 97980
rect 183520 97940 399484 97968
rect 183520 97928 183526 97940
rect 399478 97928 399484 97940
rect 399536 97928 399542 97980
rect 100754 97248 100760 97300
rect 100812 97288 100818 97300
rect 109770 97288 109776 97300
rect 100812 97260 109776 97288
rect 100812 97248 100818 97260
rect 109770 97248 109776 97260
rect 109828 97248 109834 97300
rect 183186 96568 183192 96620
rect 183244 96608 183250 96620
rect 418798 96608 418804 96620
rect 183244 96580 418804 96608
rect 183244 96568 183250 96580
rect 418798 96568 418804 96580
rect 418856 96568 418862 96620
rect 183278 95140 183284 95192
rect 183336 95180 183342 95192
rect 417418 95180 417424 95192
rect 183336 95152 417424 95180
rect 183336 95140 183342 95152
rect 417418 95140 417424 95152
rect 417476 95140 417482 95192
rect 183278 93780 183284 93832
rect 183336 93820 183342 93832
rect 414658 93820 414664 93832
rect 183336 93792 414664 93820
rect 183336 93780 183342 93792
rect 414658 93780 414664 93792
rect 414716 93780 414722 93832
rect 109770 93576 109776 93628
rect 109828 93616 109834 93628
rect 113818 93616 113824 93628
rect 109828 93588 113824 93616
rect 109828 93576 109834 93588
rect 113818 93576 113824 93588
rect 113876 93576 113882 93628
rect 109678 93236 109684 93288
rect 109736 93276 109742 93288
rect 110414 93276 110420 93288
rect 109736 93248 110420 93276
rect 109736 93236 109742 93248
rect 110414 93236 110420 93248
rect 110472 93236 110478 93288
rect 183462 92420 183468 92472
rect 183520 92460 183526 92472
rect 413278 92460 413284 92472
rect 183520 92432 413284 92460
rect 183520 92420 183526 92432
rect 413278 92420 413284 92432
rect 413336 92420 413342 92472
rect 110414 91060 110420 91112
rect 110472 91100 110478 91112
rect 110472 91072 113174 91100
rect 110472 91060 110478 91072
rect 113146 91032 113174 91072
rect 115290 91032 115296 91044
rect 113146 91004 115296 91032
rect 115290 90992 115296 91004
rect 115348 90992 115354 91044
rect 183462 89632 183468 89684
rect 183520 89672 183526 89684
rect 189718 89672 189724 89684
rect 183520 89644 189724 89672
rect 183520 89632 183526 89644
rect 189718 89632 189724 89644
rect 189776 89632 189782 89684
rect 183462 88204 183468 88256
rect 183520 88244 183526 88256
rect 188338 88244 188344 88256
rect 183520 88216 188344 88244
rect 183520 88204 183526 88216
rect 188338 88204 188344 88216
rect 188396 88204 188402 88256
rect 3142 85552 3148 85604
rect 3200 85592 3206 85604
rect 3510 85592 3516 85604
rect 3200 85564 3516 85592
rect 3200 85552 3206 85564
rect 3510 85552 3516 85564
rect 3568 85552 3574 85604
rect 3602 85552 3608 85604
rect 3660 85552 3666 85604
rect 183462 85552 183468 85604
rect 183520 85592 183526 85604
rect 580166 85592 580172 85604
rect 183520 85564 580172 85592
rect 183520 85552 183526 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 3620 85400 3648 85552
rect 3602 85348 3608 85400
rect 3660 85348 3666 85400
rect 3878 84940 3884 84992
rect 3936 84940 3942 84992
rect 3050 84804 3056 84856
rect 3108 84844 3114 84856
rect 3326 84844 3332 84856
rect 3108 84816 3332 84844
rect 3108 84804 3114 84816
rect 3326 84804 3332 84816
rect 3384 84804 3390 84856
rect 3896 84720 3924 84940
rect 3878 84668 3884 84720
rect 3936 84668 3942 84720
rect 3970 84192 3976 84244
rect 4028 84232 4034 84244
rect 120442 84232 120448 84244
rect 4028 84204 120448 84232
rect 4028 84192 4034 84204
rect 120442 84192 120448 84204
rect 120500 84192 120506 84244
rect 178954 82084 178960 82136
rect 179012 82124 179018 82136
rect 580350 82124 580356 82136
rect 179012 82096 580356 82124
rect 179012 82084 179018 82096
rect 580350 82084 580356 82096
rect 580408 82084 580414 82136
rect 183462 81404 183468 81456
rect 183520 81444 183526 81456
rect 555418 81444 555424 81456
rect 183520 81416 555424 81444
rect 183520 81404 183526 81416
rect 555418 81404 555424 81416
rect 555476 81404 555482 81456
rect 147646 80804 168788 80832
rect 113818 80656 113824 80708
rect 113876 80696 113882 80708
rect 147646 80696 147674 80804
rect 113876 80668 147674 80696
rect 153166 80736 164234 80764
rect 113876 80656 113882 80668
rect 120046 80328 142108 80356
rect 119338 79976 119344 80028
rect 119396 80016 119402 80028
rect 120046 80016 120074 80328
rect 125042 80248 125048 80300
rect 125100 80288 125106 80300
rect 125100 80260 129734 80288
rect 125100 80248 125106 80260
rect 129706 80152 129734 80260
rect 129706 80124 132494 80152
rect 123662 80044 123668 80096
rect 123720 80084 123726 80096
rect 123720 80056 128446 80084
rect 123720 80044 123726 80056
rect 119396 79988 120074 80016
rect 125566 79988 126882 80016
rect 119396 79976 119402 79988
rect 124950 79908 124956 79960
rect 125008 79948 125014 79960
rect 125566 79948 125594 79988
rect 126744 79948 126750 79960
rect 125008 79920 125594 79948
rect 126440 79920 126750 79948
rect 125008 79908 125014 79920
rect 122926 79840 122932 79892
rect 122984 79880 122990 79892
rect 126008 79880 126014 79892
rect 122984 79852 126014 79880
rect 122984 79840 122990 79852
rect 126008 79840 126014 79852
rect 126066 79840 126072 79892
rect 126284 79840 126290 79892
rect 126342 79840 126348 79892
rect 125502 79772 125508 79824
rect 125560 79812 125566 79824
rect 125916 79812 125922 79824
rect 125560 79784 125922 79812
rect 125560 79772 125566 79784
rect 125916 79772 125922 79784
rect 125974 79772 125980 79824
rect 126302 79812 126330 79840
rect 126072 79784 126330 79812
rect 126072 79756 126100 79784
rect 126054 79704 126060 79756
rect 126112 79704 126118 79756
rect 126330 79704 126336 79756
rect 126388 79744 126394 79756
rect 126440 79744 126468 79920
rect 126744 79908 126750 79920
rect 126802 79908 126808 79960
rect 126560 79840 126566 79892
rect 126618 79840 126624 79892
rect 126652 79840 126658 79892
rect 126710 79880 126716 79892
rect 126854 79880 126882 79988
rect 128418 79960 128446 80056
rect 126928 79908 126934 79960
rect 126986 79908 126992 79960
rect 127020 79908 127026 79960
rect 127078 79908 127084 79960
rect 127480 79908 127486 79960
rect 127538 79908 127544 79960
rect 127756 79908 127762 79960
rect 127814 79908 127820 79960
rect 128032 79908 128038 79960
rect 128090 79908 128096 79960
rect 128216 79908 128222 79960
rect 128274 79908 128280 79960
rect 128400 79908 128406 79960
rect 128458 79908 128464 79960
rect 129044 79948 129050 79960
rect 128786 79920 129050 79948
rect 126710 79852 126882 79880
rect 126710 79840 126716 79852
rect 126578 79812 126606 79840
rect 126946 79812 126974 79908
rect 126388 79716 126468 79744
rect 126532 79784 126606 79812
rect 126808 79784 126974 79812
rect 127038 79824 127066 79908
rect 127038 79784 127072 79824
rect 126388 79704 126394 79716
rect 5166 79568 5172 79620
rect 5224 79608 5230 79620
rect 120718 79608 120724 79620
rect 5224 79580 120724 79608
rect 5224 79568 5230 79580
rect 120718 79568 120724 79580
rect 120776 79568 120782 79620
rect 126532 79608 126560 79784
rect 125888 79580 126560 79608
rect 125888 79552 125916 79580
rect 115906 79512 120074 79540
rect 115198 79432 115204 79484
rect 115256 79472 115262 79484
rect 115906 79472 115934 79512
rect 115256 79444 115934 79472
rect 120046 79472 120074 79512
rect 125870 79500 125876 79552
rect 125928 79500 125934 79552
rect 125962 79500 125968 79552
rect 126020 79540 126026 79552
rect 126808 79540 126836 79784
rect 127066 79772 127072 79784
rect 127124 79772 127130 79824
rect 126974 79704 126980 79756
rect 127032 79744 127038 79756
rect 127498 79744 127526 79908
rect 127664 79840 127670 79892
rect 127722 79840 127728 79892
rect 127032 79716 127526 79744
rect 127032 79704 127038 79716
rect 126882 79636 126888 79688
rect 126940 79676 126946 79688
rect 127682 79676 127710 79840
rect 126940 79648 127710 79676
rect 126940 79636 126946 79648
rect 126020 79512 126836 79540
rect 126020 79500 126026 79512
rect 127158 79500 127164 79552
rect 127216 79540 127222 79552
rect 127774 79540 127802 79908
rect 128050 79824 128078 79908
rect 128234 79824 128262 79908
rect 128050 79784 128084 79824
rect 128078 79772 128084 79784
rect 128136 79772 128142 79824
rect 128170 79772 128176 79824
rect 128228 79784 128262 79824
rect 128228 79772 128234 79784
rect 128354 79568 128360 79620
rect 128412 79608 128418 79620
rect 128786 79608 128814 79920
rect 129044 79908 129050 79920
rect 129102 79908 129108 79960
rect 129136 79908 129142 79960
rect 129194 79908 129200 79960
rect 129320 79908 129326 79960
rect 129378 79908 129384 79960
rect 129596 79908 129602 79960
rect 129654 79908 129660 79960
rect 129688 79908 129694 79960
rect 129746 79908 129752 79960
rect 129780 79908 129786 79960
rect 129838 79908 129844 79960
rect 129964 79908 129970 79960
rect 130022 79948 130028 79960
rect 130022 79920 130378 79948
rect 130022 79908 130028 79920
rect 128952 79880 128958 79892
rect 128924 79840 128958 79880
rect 129010 79840 129016 79892
rect 128924 79756 128952 79840
rect 129154 79756 129182 79908
rect 129338 79812 129366 79908
rect 129412 79840 129418 79892
rect 129470 79840 129476 79892
rect 129504 79840 129510 79892
rect 129562 79840 129568 79892
rect 128906 79704 128912 79756
rect 128964 79704 128970 79756
rect 129090 79704 129096 79756
rect 129148 79716 129182 79756
rect 129292 79784 129366 79812
rect 129148 79704 129154 79716
rect 129292 79688 129320 79784
rect 129430 79744 129458 79840
rect 129384 79716 129458 79744
rect 129384 79688 129412 79716
rect 129274 79636 129280 79688
rect 129332 79636 129338 79688
rect 129366 79636 129372 79688
rect 129424 79636 129430 79688
rect 129522 79676 129550 79840
rect 129476 79648 129550 79676
rect 129476 79620 129504 79648
rect 129614 79620 129642 79908
rect 129706 79744 129734 79908
rect 129798 79824 129826 79908
rect 130148 79880 130154 79892
rect 130120 79840 130154 79880
rect 130206 79840 130212 79892
rect 130240 79840 130246 79892
rect 130298 79840 130304 79892
rect 129780 79772 129786 79824
rect 129838 79772 129844 79824
rect 129706 79716 129872 79744
rect 129844 79688 129872 79716
rect 129826 79636 129832 79688
rect 129884 79636 129890 79688
rect 129918 79636 129924 79688
rect 129976 79676 129982 79688
rect 130120 79676 130148 79840
rect 130258 79756 130286 79840
rect 130194 79704 130200 79756
rect 130252 79716 130286 79756
rect 130252 79704 130258 79716
rect 130350 79676 130378 79920
rect 130516 79908 130522 79960
rect 130574 79908 130580 79960
rect 130976 79948 130982 79960
rect 130626 79920 130982 79948
rect 130534 79688 130562 79908
rect 129976 79648 130148 79676
rect 130212 79648 130378 79676
rect 129976 79636 129982 79648
rect 128412 79580 128814 79608
rect 128412 79568 128418 79580
rect 129458 79568 129464 79620
rect 129516 79568 129522 79620
rect 129550 79568 129556 79620
rect 129608 79580 129642 79620
rect 129608 79568 129614 79580
rect 130010 79568 130016 79620
rect 130068 79608 130074 79620
rect 130212 79608 130240 79648
rect 130470 79636 130476 79688
rect 130528 79648 130562 79688
rect 130528 79636 130534 79648
rect 130068 79580 130240 79608
rect 130068 79568 130074 79580
rect 127216 79512 127802 79540
rect 127216 79500 127222 79512
rect 128538 79500 128544 79552
rect 128596 79540 128602 79552
rect 130626 79540 130654 79920
rect 130976 79908 130982 79920
rect 131034 79908 131040 79960
rect 131528 79908 131534 79960
rect 131586 79908 131592 79960
rect 131712 79908 131718 79960
rect 131770 79908 131776 79960
rect 130884 79840 130890 79892
rect 130942 79840 130948 79892
rect 131160 79880 131166 79892
rect 131040 79852 131166 79880
rect 130902 79756 130930 79840
rect 130902 79716 130936 79756
rect 130930 79704 130936 79716
rect 130988 79704 130994 79756
rect 131040 79552 131068 79852
rect 131160 79840 131166 79852
rect 131218 79840 131224 79892
rect 131344 79840 131350 79892
rect 131402 79840 131408 79892
rect 131206 79636 131212 79688
rect 131264 79676 131270 79688
rect 131362 79676 131390 79840
rect 131546 79824 131574 79908
rect 131482 79772 131488 79824
rect 131540 79784 131574 79824
rect 131540 79772 131546 79784
rect 131730 79756 131758 79908
rect 132466 79892 132494 80124
rect 137710 79988 138842 80016
rect 137710 79960 137738 79988
rect 132908 79948 132914 79960
rect 132650 79920 132914 79948
rect 131988 79840 131994 79892
rect 132046 79840 132052 79892
rect 132264 79840 132270 79892
rect 132322 79840 132328 79892
rect 132448 79840 132454 79892
rect 132506 79840 132512 79892
rect 131804 79772 131810 79824
rect 131862 79772 131868 79824
rect 131666 79704 131672 79756
rect 131724 79716 131758 79756
rect 131724 79704 131730 79716
rect 131822 79688 131850 79772
rect 131264 79648 131390 79676
rect 131264 79636 131270 79648
rect 131758 79636 131764 79688
rect 131816 79648 131850 79688
rect 131816 79636 131822 79648
rect 132006 79552 132034 79840
rect 128596 79512 130654 79540
rect 128596 79500 128602 79512
rect 131022 79500 131028 79552
rect 131080 79500 131086 79552
rect 132006 79512 132040 79552
rect 132034 79500 132040 79512
rect 132092 79500 132098 79552
rect 132282 79540 132310 79840
rect 132540 79772 132546 79824
rect 132598 79772 132604 79824
rect 132402 79636 132408 79688
rect 132460 79676 132466 79688
rect 132558 79676 132586 79772
rect 132460 79648 132586 79676
rect 132460 79636 132466 79648
rect 132650 79620 132678 79920
rect 132908 79908 132914 79920
rect 132966 79908 132972 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134288 79908 134294 79960
rect 134346 79908 134352 79960
rect 135024 79948 135030 79960
rect 134996 79908 135030 79948
rect 135082 79908 135088 79960
rect 135116 79908 135122 79960
rect 135174 79908 135180 79960
rect 135484 79908 135490 79960
rect 135542 79908 135548 79960
rect 136588 79948 136594 79960
rect 136008 79920 136594 79948
rect 132816 79840 132822 79892
rect 132874 79840 132880 79892
rect 133184 79840 133190 79892
rect 133242 79840 133248 79892
rect 133736 79840 133742 79892
rect 133794 79840 133800 79892
rect 132586 79568 132592 79620
rect 132644 79580 132678 79620
rect 132644 79568 132650 79580
rect 132834 79552 132862 79840
rect 132678 79540 132684 79552
rect 132282 79512 132684 79540
rect 132678 79500 132684 79512
rect 132736 79500 132742 79552
rect 132770 79500 132776 79552
rect 132828 79512 132862 79552
rect 132828 79500 132834 79512
rect 133046 79500 133052 79552
rect 133104 79540 133110 79552
rect 133202 79540 133230 79840
rect 133368 79812 133374 79824
rect 133340 79772 133374 79812
rect 133426 79772 133432 79824
rect 133644 79772 133650 79824
rect 133702 79772 133708 79824
rect 133340 79552 133368 79772
rect 133662 79620 133690 79772
rect 133598 79568 133604 79620
rect 133656 79580 133690 79620
rect 133656 79568 133662 79580
rect 133754 79552 133782 79840
rect 133938 79824 133966 79908
rect 133874 79772 133880 79824
rect 133932 79784 133966 79824
rect 133932 79772 133938 79784
rect 134122 79688 134150 79908
rect 134058 79636 134064 79688
rect 134116 79648 134150 79688
rect 134116 79636 134122 79648
rect 134150 79568 134156 79620
rect 134208 79608 134214 79620
rect 134306 79608 134334 79908
rect 134564 79840 134570 79892
rect 134622 79840 134628 79892
rect 134748 79840 134754 79892
rect 134806 79880 134812 79892
rect 134806 79840 134840 79880
rect 134208 79580 134334 79608
rect 134208 79568 134214 79580
rect 134426 79568 134432 79620
rect 134484 79608 134490 79620
rect 134582 79608 134610 79840
rect 134484 79580 134610 79608
rect 134484 79568 134490 79580
rect 133104 79512 133230 79540
rect 133104 79500 133110 79512
rect 133322 79500 133328 79552
rect 133380 79500 133386 79552
rect 133690 79500 133696 79552
rect 133748 79512 133782 79552
rect 133748 79500 133754 79512
rect 133966 79500 133972 79552
rect 134024 79540 134030 79552
rect 134812 79540 134840 79840
rect 134996 79620 135024 79908
rect 135134 79880 135162 79908
rect 135088 79852 135162 79880
rect 135088 79620 135116 79852
rect 135300 79812 135306 79824
rect 135180 79784 135306 79812
rect 134978 79568 134984 79620
rect 135036 79568 135042 79620
rect 135070 79568 135076 79620
rect 135128 79568 135134 79620
rect 134024 79512 134840 79540
rect 134024 79500 134030 79512
rect 134058 79472 134064 79484
rect 120046 79444 134064 79472
rect 115256 79432 115262 79444
rect 134058 79432 134064 79444
rect 134116 79432 134122 79484
rect 120718 79364 120724 79416
rect 120776 79404 120782 79416
rect 120776 79376 133874 79404
rect 120776 79364 120782 79376
rect 125318 79296 125324 79348
rect 125376 79336 125382 79348
rect 126238 79336 126244 79348
rect 125376 79308 126244 79336
rect 125376 79296 125382 79308
rect 126238 79296 126244 79308
rect 126296 79296 126302 79348
rect 133846 79268 133874 79376
rect 134518 79296 134524 79348
rect 134576 79336 134582 79348
rect 135180 79336 135208 79784
rect 135300 79772 135306 79784
rect 135358 79772 135364 79824
rect 135502 79552 135530 79908
rect 135668 79880 135674 79892
rect 135640 79840 135674 79880
rect 135726 79840 135732 79892
rect 135640 79688 135668 79840
rect 135622 79636 135628 79688
rect 135680 79636 135686 79688
rect 136008 79552 136036 79920
rect 136588 79908 136594 79920
rect 136646 79908 136652 79960
rect 137416 79948 137422 79960
rect 137388 79908 137422 79948
rect 137474 79908 137480 79960
rect 137508 79908 137514 79960
rect 137566 79908 137572 79960
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137692 79908 137698 79960
rect 137750 79908 137756 79960
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138520 79948 138526 79960
rect 138492 79908 138526 79948
rect 138578 79908 138584 79960
rect 138612 79908 138618 79960
rect 138670 79908 138676 79960
rect 136128 79840 136134 79892
rect 136186 79840 136192 79892
rect 136312 79840 136318 79892
rect 136370 79840 136376 79892
rect 136404 79840 136410 79892
rect 136462 79840 136468 79892
rect 136956 79840 136962 79892
rect 137014 79840 137020 79892
rect 137048 79840 137054 79892
rect 137106 79880 137112 79892
rect 137106 79840 137140 79880
rect 137232 79840 137238 79892
rect 137290 79880 137296 79892
rect 137290 79840 137324 79880
rect 135502 79512 135536 79552
rect 135530 79500 135536 79512
rect 135588 79500 135594 79552
rect 135990 79500 135996 79552
rect 136048 79500 136054 79552
rect 135346 79364 135352 79416
rect 135404 79404 135410 79416
rect 136146 79404 136174 79840
rect 136330 79608 136358 79840
rect 136284 79580 136358 79608
rect 136284 79552 136312 79580
rect 136422 79552 136450 79840
rect 136496 79772 136502 79824
rect 136554 79772 136560 79824
rect 136772 79812 136778 79824
rect 136744 79772 136778 79812
rect 136830 79772 136836 79824
rect 136864 79772 136870 79824
rect 136922 79772 136928 79824
rect 136514 79620 136542 79772
rect 136744 79688 136772 79772
rect 136726 79636 136732 79688
rect 136784 79636 136790 79688
rect 136882 79676 136910 79772
rect 136836 79648 136910 79676
rect 136514 79580 136548 79620
rect 136542 79568 136548 79580
rect 136600 79568 136606 79620
rect 136266 79500 136272 79552
rect 136324 79500 136330 79552
rect 136358 79500 136364 79552
rect 136416 79512 136450 79552
rect 136836 79540 136864 79648
rect 136974 79620 137002 79840
rect 137112 79756 137140 79840
rect 137296 79756 137324 79840
rect 137094 79704 137100 79756
rect 137152 79704 137158 79756
rect 137278 79704 137284 79756
rect 137336 79704 137342 79756
rect 137388 79688 137416 79908
rect 137370 79636 137376 79688
rect 137428 79636 137434 79688
rect 136910 79568 136916 79620
rect 136968 79580 137002 79620
rect 136968 79568 136974 79580
rect 137526 79552 137554 79908
rect 137002 79540 137008 79552
rect 136836 79512 137008 79540
rect 136416 79500 136422 79512
rect 137002 79500 137008 79512
rect 137060 79500 137066 79552
rect 137462 79500 137468 79552
rect 137520 79512 137554 79552
rect 137520 79500 137526 79512
rect 136726 79432 136732 79484
rect 136784 79472 136790 79484
rect 137618 79472 137646 79908
rect 138078 79688 138106 79908
rect 138152 79840 138158 79892
rect 138210 79840 138216 79892
rect 138244 79840 138250 79892
rect 138302 79840 138308 79892
rect 138014 79636 138020 79688
rect 138072 79648 138106 79688
rect 138072 79636 138078 79648
rect 136784 79444 137646 79472
rect 136784 79432 136790 79444
rect 135404 79376 136174 79404
rect 135404 79364 135410 79376
rect 134576 79308 135208 79336
rect 138170 79336 138198 79840
rect 138262 79540 138290 79840
rect 138492 79620 138520 79908
rect 138630 79880 138658 79908
rect 138814 79880 138842 79988
rect 141298 79988 141786 80016
rect 141298 79960 141326 79988
rect 139256 79908 139262 79960
rect 139314 79908 139320 79960
rect 139348 79908 139354 79960
rect 139406 79908 139412 79960
rect 139440 79908 139446 79960
rect 139498 79908 139504 79960
rect 139808 79948 139814 79960
rect 139550 79920 139814 79948
rect 138584 79852 138658 79880
rect 138768 79852 138842 79880
rect 138474 79568 138480 79620
rect 138532 79568 138538 79620
rect 138382 79540 138388 79552
rect 138262 79512 138388 79540
rect 138382 79500 138388 79512
rect 138440 79500 138446 79552
rect 138584 79472 138612 79852
rect 138768 79620 138796 79852
rect 138888 79840 138894 79892
rect 138946 79880 138952 79892
rect 138946 79840 138980 79880
rect 138750 79568 138756 79620
rect 138808 79568 138814 79620
rect 138952 79608 138980 79840
rect 139072 79772 139078 79824
rect 139130 79812 139136 79824
rect 139130 79772 139164 79812
rect 139136 79620 139164 79772
rect 139026 79608 139032 79620
rect 138952 79580 139032 79608
rect 139026 79568 139032 79580
rect 139084 79568 139090 79620
rect 139118 79568 139124 79620
rect 139176 79568 139182 79620
rect 138934 79472 138940 79484
rect 138584 79444 138940 79472
rect 138934 79432 138940 79444
rect 138992 79432 138998 79484
rect 139274 79404 139302 79908
rect 139366 79472 139394 79908
rect 139458 79824 139486 79908
rect 139440 79772 139446 79824
rect 139498 79772 139504 79824
rect 139550 79688 139578 79920
rect 139808 79908 139814 79920
rect 139866 79908 139872 79960
rect 140084 79908 140090 79960
rect 140142 79908 140148 79960
rect 140268 79948 140274 79960
rect 140240 79908 140274 79948
rect 140326 79908 140332 79960
rect 140360 79908 140366 79960
rect 140418 79908 140424 79960
rect 140544 79908 140550 79960
rect 140602 79908 140608 79960
rect 140728 79908 140734 79960
rect 140786 79908 140792 79960
rect 140820 79908 140826 79960
rect 140878 79908 140884 79960
rect 141188 79908 141194 79960
rect 141246 79908 141252 79960
rect 141280 79908 141286 79960
rect 141338 79908 141344 79960
rect 141372 79908 141378 79960
rect 141430 79908 141436 79960
rect 141556 79908 141562 79960
rect 141614 79908 141620 79960
rect 141648 79908 141654 79960
rect 141706 79908 141712 79960
rect 139624 79840 139630 79892
rect 139682 79840 139688 79892
rect 139900 79880 139906 79892
rect 139872 79840 139906 79880
rect 139958 79840 139964 79892
rect 139486 79636 139492 79688
rect 139544 79648 139578 79688
rect 139544 79636 139550 79648
rect 139642 79540 139670 79840
rect 139872 79756 139900 79840
rect 139854 79704 139860 79756
rect 139912 79704 139918 79756
rect 139946 79704 139952 79756
rect 140004 79744 140010 79756
rect 140102 79744 140130 79908
rect 140004 79716 140130 79744
rect 140004 79704 140010 79716
rect 140240 79620 140268 79908
rect 140378 79880 140406 79908
rect 140332 79852 140406 79880
rect 140332 79824 140360 79852
rect 140314 79772 140320 79824
rect 140372 79772 140378 79824
rect 140562 79688 140590 79908
rect 140746 79812 140774 79908
rect 140700 79784 140774 79812
rect 140700 79756 140728 79784
rect 140838 79756 140866 79908
rect 140912 79840 140918 79892
rect 140970 79840 140976 79892
rect 141004 79840 141010 79892
rect 141062 79840 141068 79892
rect 140682 79704 140688 79756
rect 140740 79704 140746 79756
rect 140774 79704 140780 79756
rect 140832 79716 140866 79756
rect 140832 79704 140838 79716
rect 140562 79648 140596 79688
rect 140590 79636 140596 79648
rect 140648 79636 140654 79688
rect 140930 79620 140958 79840
rect 141022 79812 141050 79840
rect 141022 79784 141096 79812
rect 141068 79620 141096 79784
rect 140222 79568 140228 79620
rect 140280 79568 140286 79620
rect 140866 79568 140872 79620
rect 140924 79580 140958 79620
rect 140924 79568 140930 79580
rect 141050 79568 141056 79620
rect 141108 79568 141114 79620
rect 139762 79540 139768 79552
rect 139642 79512 139768 79540
rect 139762 79500 139768 79512
rect 139820 79500 139826 79552
rect 140958 79500 140964 79552
rect 141016 79540 141022 79552
rect 141206 79540 141234 79908
rect 141390 79812 141418 79908
rect 141464 79840 141470 79892
rect 141522 79840 141528 79892
rect 141016 79512 141234 79540
rect 141344 79784 141418 79812
rect 141016 79500 141022 79512
rect 139946 79472 139952 79484
rect 139366 79444 139952 79472
rect 139946 79432 139952 79444
rect 140004 79432 140010 79484
rect 141344 79416 141372 79784
rect 141482 79744 141510 79840
rect 141436 79716 141510 79744
rect 141436 79416 141464 79716
rect 141574 79676 141602 79908
rect 141528 79648 141602 79676
rect 141528 79552 141556 79648
rect 141666 79620 141694 79908
rect 141602 79568 141608 79620
rect 141660 79580 141694 79620
rect 141660 79568 141666 79580
rect 141758 79552 141786 79988
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 141510 79500 141516 79552
rect 141568 79500 141574 79552
rect 141694 79500 141700 79552
rect 141752 79512 141786 79552
rect 141752 79500 141758 79512
rect 141942 79416 141970 79908
rect 142080 79552 142108 80328
rect 149118 80260 153102 80288
rect 142402 80056 144868 80084
rect 142402 79960 142430 80056
rect 142678 79988 143442 80016
rect 142678 79960 142706 79988
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 142384 79908 142390 79960
rect 142442 79908 142448 79960
rect 142476 79908 142482 79960
rect 142534 79908 142540 79960
rect 142568 79908 142574 79960
rect 142626 79908 142632 79960
rect 142660 79908 142666 79960
rect 142718 79908 142724 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 142218 79620 142246 79908
rect 142494 79812 142522 79908
rect 142586 79880 142614 79908
rect 142586 79852 142844 79880
rect 142706 79812 142712 79824
rect 142494 79784 142712 79812
rect 142706 79772 142712 79784
rect 142764 79772 142770 79824
rect 142816 79688 142844 79852
rect 142936 79772 142942 79824
rect 142994 79772 143000 79824
rect 143028 79772 143034 79824
rect 143086 79772 143092 79824
rect 143120 79772 143126 79824
rect 143178 79772 143184 79824
rect 143230 79812 143258 79908
rect 143230 79784 143304 79812
rect 142954 79744 142982 79772
rect 142908 79716 142982 79744
rect 142798 79636 142804 79688
rect 142856 79636 142862 79688
rect 142218 79580 142252 79620
rect 142246 79568 142252 79580
rect 142304 79568 142310 79620
rect 142062 79500 142068 79552
rect 142120 79500 142126 79552
rect 142908 79540 142936 79716
rect 143046 79688 143074 79772
rect 143138 79744 143166 79772
rect 143138 79716 143212 79744
rect 143184 79688 143212 79716
rect 143276 79688 143304 79784
rect 142982 79636 142988 79688
rect 143040 79648 143074 79688
rect 143040 79636 143046 79648
rect 143166 79636 143172 79688
rect 143224 79636 143230 79688
rect 143258 79636 143264 79688
rect 143316 79636 143322 79688
rect 143074 79568 143080 79620
rect 143132 79608 143138 79620
rect 143414 79608 143442 79988
rect 143764 79908 143770 79960
rect 143822 79908 143828 79960
rect 143856 79908 143862 79960
rect 143914 79948 143920 79960
rect 143914 79920 144316 79948
rect 143914 79908 143920 79920
rect 143132 79580 143442 79608
rect 143782 79608 143810 79908
rect 144132 79840 144138 79892
rect 144190 79880 144196 79892
rect 144190 79840 144224 79880
rect 144040 79772 144046 79824
rect 144098 79772 144104 79824
rect 144058 79744 144086 79772
rect 144058 79716 144132 79744
rect 144104 79620 144132 79716
rect 144196 79620 144224 79840
rect 144288 79620 144316 79920
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144500 79908 144506 79960
rect 144558 79908 144564 79960
rect 144684 79908 144690 79960
rect 144742 79908 144748 79960
rect 143902 79608 143908 79620
rect 143782 79580 143908 79608
rect 143132 79568 143138 79580
rect 143902 79568 143908 79580
rect 143960 79568 143966 79620
rect 144086 79568 144092 79620
rect 144144 79568 144150 79620
rect 144178 79568 144184 79620
rect 144236 79568 144242 79620
rect 144270 79568 144276 79620
rect 144328 79568 144334 79620
rect 143442 79540 143448 79552
rect 142908 79512 143448 79540
rect 143442 79500 143448 79512
rect 143500 79500 143506 79552
rect 143534 79500 143540 79552
rect 143592 79540 143598 79552
rect 144426 79540 144454 79908
rect 144518 79756 144546 79908
rect 144702 79756 144730 79908
rect 144518 79716 144552 79756
rect 144546 79704 144552 79716
rect 144604 79704 144610 79756
rect 144638 79704 144644 79756
rect 144696 79716 144730 79756
rect 144696 79704 144702 79716
rect 144840 79620 144868 80056
rect 145070 79988 145466 80016
rect 144960 79772 144966 79824
rect 145018 79772 145024 79824
rect 144978 79744 145006 79772
rect 144932 79716 145006 79744
rect 144932 79688 144960 79716
rect 145070 79688 145098 79988
rect 145438 79960 145466 79988
rect 149118 79960 149146 80260
rect 150360 79988 150802 80016
rect 145144 79908 145150 79960
rect 145202 79908 145208 79960
rect 145420 79908 145426 79960
rect 145478 79908 145484 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 145880 79908 145886 79960
rect 145938 79948 145944 79960
rect 145938 79920 146018 79948
rect 145938 79908 145944 79920
rect 144914 79636 144920 79688
rect 144972 79636 144978 79688
rect 145006 79636 145012 79688
rect 145064 79648 145098 79688
rect 145064 79636 145070 79648
rect 144822 79568 144828 79620
rect 144880 79568 144886 79620
rect 143592 79512 144454 79540
rect 145162 79540 145190 79908
rect 145604 79840 145610 79892
rect 145662 79840 145668 79892
rect 145622 79688 145650 79840
rect 145806 79824 145834 79908
rect 145806 79784 145840 79824
rect 145834 79772 145840 79784
rect 145892 79772 145898 79824
rect 145622 79648 145656 79688
rect 145650 79636 145656 79648
rect 145708 79636 145714 79688
rect 145990 79552 146018 79920
rect 147076 79908 147082 79960
rect 147134 79908 147140 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 148088 79908 148094 79960
rect 148146 79908 148152 79960
rect 148180 79908 148186 79960
rect 148238 79908 148244 79960
rect 148272 79908 148278 79960
rect 148330 79908 148336 79960
rect 149008 79908 149014 79960
rect 149066 79908 149072 79960
rect 149100 79908 149106 79960
rect 149158 79908 149164 79960
rect 149468 79948 149474 79960
rect 149256 79920 149474 79948
rect 146984 79840 146990 79892
rect 147042 79840 147048 79892
rect 146616 79772 146622 79824
rect 146674 79772 146680 79824
rect 146634 79608 146662 79772
rect 146312 79580 146662 79608
rect 147002 79608 147030 79840
rect 147094 79688 147122 79908
rect 147260 79840 147266 79892
rect 147318 79840 147324 79892
rect 147278 79744 147306 79840
rect 147462 79824 147490 79908
rect 147904 79840 147910 79892
rect 147962 79840 147968 79892
rect 147398 79772 147404 79824
rect 147456 79784 147490 79824
rect 147456 79772 147462 79784
rect 147720 79772 147726 79824
rect 147778 79772 147784 79824
rect 147812 79772 147818 79824
rect 147870 79772 147876 79824
rect 147278 79716 147536 79744
rect 147094 79648 147128 79688
rect 147122 79636 147128 79648
rect 147180 79636 147186 79688
rect 147214 79608 147220 79620
rect 147002 79580 147220 79608
rect 146312 79552 146340 79580
rect 147214 79568 147220 79580
rect 147272 79568 147278 79620
rect 147508 79552 147536 79716
rect 147738 79620 147766 79772
rect 147830 79688 147858 79772
rect 147922 79756 147950 79840
rect 148106 79756 148134 79908
rect 147922 79716 147956 79756
rect 147950 79704 147956 79716
rect 148008 79704 148014 79756
rect 148042 79704 148048 79756
rect 148100 79716 148134 79756
rect 148100 79704 148106 79716
rect 147830 79648 147864 79688
rect 147858 79636 147864 79648
rect 147916 79636 147922 79688
rect 147738 79580 147772 79620
rect 147766 79568 147772 79580
rect 147824 79568 147830 79620
rect 145374 79540 145380 79552
rect 145162 79512 145380 79540
rect 143592 79500 143598 79512
rect 145374 79500 145380 79512
rect 145432 79500 145438 79552
rect 145990 79512 146024 79552
rect 146018 79500 146024 79512
rect 146076 79500 146082 79552
rect 146294 79500 146300 79552
rect 146352 79500 146358 79552
rect 147490 79500 147496 79552
rect 147548 79500 147554 79552
rect 148198 79540 148226 79908
rect 148290 79824 148318 79908
rect 148364 79840 148370 79892
rect 148422 79840 148428 79892
rect 148824 79840 148830 79892
rect 148882 79840 148888 79892
rect 148272 79772 148278 79824
rect 148330 79772 148336 79824
rect 148382 79688 148410 79840
rect 148842 79756 148870 79840
rect 148778 79704 148784 79756
rect 148836 79716 148870 79756
rect 148836 79704 148842 79716
rect 148318 79636 148324 79688
rect 148376 79648 148410 79688
rect 149026 79688 149054 79908
rect 149256 79688 149284 79920
rect 149468 79908 149474 79920
rect 149526 79908 149532 79960
rect 149744 79908 149750 79960
rect 149802 79948 149808 79960
rect 149802 79920 149928 79948
rect 149802 79908 149808 79920
rect 149376 79840 149382 79892
rect 149434 79880 149440 79892
rect 149434 79852 149836 79880
rect 149434 79840 149440 79852
rect 149808 79688 149836 79852
rect 149026 79648 149060 79688
rect 148376 79636 148382 79648
rect 149054 79636 149060 79648
rect 149112 79636 149118 79688
rect 149238 79636 149244 79688
rect 149296 79636 149302 79688
rect 149790 79636 149796 79688
rect 149848 79636 149854 79688
rect 149900 79620 149928 79920
rect 150020 79908 150026 79960
rect 150078 79908 150084 79960
rect 148870 79568 148876 79620
rect 148928 79608 148934 79620
rect 148928 79580 149698 79608
rect 148928 79568 148934 79580
rect 149514 79540 149520 79552
rect 148198 79512 149520 79540
rect 149514 79500 149520 79512
rect 149572 79500 149578 79552
rect 149670 79540 149698 79580
rect 149882 79568 149888 79620
rect 149940 79568 149946 79620
rect 150038 79540 150066 79908
rect 150112 79840 150118 79892
rect 150170 79840 150176 79892
rect 150130 79756 150158 79840
rect 150130 79716 150164 79756
rect 150158 79704 150164 79716
rect 150216 79704 150222 79756
rect 150360 79620 150388 79988
rect 150774 79960 150802 79988
rect 150480 79908 150486 79960
rect 150538 79908 150544 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 151216 79908 151222 79960
rect 151274 79908 151280 79960
rect 151492 79908 151498 79960
rect 151550 79908 151556 79960
rect 151584 79908 151590 79960
rect 151642 79908 151648 79960
rect 151676 79908 151682 79960
rect 151734 79908 151740 79960
rect 151952 79948 151958 79960
rect 151786 79920 151958 79948
rect 150498 79744 150526 79908
rect 151234 79880 151262 79908
rect 150452 79716 150526 79744
rect 150820 79852 151262 79880
rect 150342 79568 150348 79620
rect 150400 79568 150406 79620
rect 149670 79512 150066 79540
rect 150452 79540 150480 79716
rect 150820 79688 150848 79852
rect 150940 79812 150946 79824
rect 150912 79772 150946 79812
rect 150998 79772 151004 79824
rect 150912 79688 150940 79772
rect 150802 79636 150808 79688
rect 150860 79636 150866 79688
rect 150894 79636 150900 79688
rect 150952 79636 150958 79688
rect 150986 79636 150992 79688
rect 151044 79676 151050 79688
rect 151510 79676 151538 79908
rect 151044 79648 151538 79676
rect 151044 79636 151050 79648
rect 151170 79568 151176 79620
rect 151228 79608 151234 79620
rect 151602 79608 151630 79908
rect 151228 79580 151630 79608
rect 151228 79568 151234 79580
rect 151694 79552 151722 79908
rect 151786 79756 151814 79920
rect 151952 79908 151958 79920
rect 152010 79908 152016 79960
rect 152044 79908 152050 79960
rect 152102 79908 152108 79960
rect 152136 79908 152142 79960
rect 152194 79908 152200 79960
rect 152504 79908 152510 79960
rect 152562 79908 152568 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 151860 79840 151866 79892
rect 151918 79880 151924 79892
rect 151918 79840 151952 79880
rect 151786 79716 151820 79756
rect 151814 79704 151820 79716
rect 151872 79704 151878 79756
rect 151924 79620 151952 79840
rect 151906 79568 151912 79620
rect 151964 79568 151970 79620
rect 151538 79540 151544 79552
rect 150452 79512 151544 79540
rect 151538 79500 151544 79512
rect 151596 79500 151602 79552
rect 151694 79512 151728 79552
rect 151722 79500 151728 79512
rect 151780 79500 151786 79552
rect 152062 79540 152090 79908
rect 152154 79608 152182 79908
rect 152522 79824 152550 79908
rect 152688 79840 152694 79892
rect 152746 79840 152752 79892
rect 152522 79784 152556 79824
rect 152550 79772 152556 79784
rect 152608 79772 152614 79824
rect 152458 79608 152464 79620
rect 152154 79580 152464 79608
rect 152458 79568 152464 79580
rect 152516 79568 152522 79620
rect 152706 79608 152734 79840
rect 152982 79688 153010 79908
rect 153074 79744 153102 80260
rect 153166 79812 153194 80736
rect 164206 80628 164234 80736
rect 168760 80696 168788 80804
rect 178494 80724 178500 80776
rect 178552 80764 178558 80776
rect 393958 80764 393964 80776
rect 178552 80736 393964 80764
rect 178552 80724 178558 80736
rect 393958 80724 393964 80736
rect 394016 80724 394022 80776
rect 174722 80696 174728 80708
rect 168760 80668 174728 80696
rect 174722 80656 174728 80668
rect 174780 80656 174786 80708
rect 504450 80696 504456 80708
rect 182146 80668 504456 80696
rect 164206 80600 168650 80628
rect 168622 80560 168650 80600
rect 174538 80560 174544 80572
rect 168622 80532 168696 80560
rect 156938 80464 162854 80492
rect 156938 80424 156966 80464
rect 153258 80396 156966 80424
rect 157030 80396 158714 80424
rect 153258 79960 153286 80396
rect 157030 80288 157058 80396
rect 156938 80260 157058 80288
rect 156938 80152 156966 80260
rect 158686 80220 158714 80396
rect 162826 80288 162854 80464
rect 168668 80424 168696 80532
rect 173038 80532 174544 80560
rect 173038 80424 173066 80532
rect 174538 80520 174544 80532
rect 174596 80520 174602 80572
rect 176010 80520 176016 80572
rect 176068 80560 176074 80572
rect 182146 80560 182174 80668
rect 504450 80656 504456 80668
rect 504508 80656 504514 80708
rect 176068 80532 182174 80560
rect 176068 80520 176074 80532
rect 176102 80492 176108 80504
rect 168668 80396 173066 80424
rect 173866 80464 176108 80492
rect 173866 80356 173894 80464
rect 176102 80452 176108 80464
rect 176160 80452 176166 80504
rect 175274 80384 175280 80436
rect 175332 80424 175338 80436
rect 182174 80424 182180 80436
rect 175332 80396 182180 80424
rect 175332 80384 175338 80396
rect 182174 80384 182180 80396
rect 182232 80384 182238 80436
rect 163424 80328 173894 80356
rect 162826 80260 163084 80288
rect 158686 80192 161474 80220
rect 154546 80124 156966 80152
rect 154546 80084 154574 80124
rect 154500 80056 154574 80084
rect 159054 80056 161382 80084
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153608 79948 153614 79960
rect 153442 79920 153614 79948
rect 153166 79784 153332 79812
rect 153074 79716 153240 79744
rect 152982 79648 153016 79688
rect 153010 79636 153016 79648
rect 153068 79636 153074 79688
rect 152918 79608 152924 79620
rect 152706 79580 152924 79608
rect 152918 79568 152924 79580
rect 152976 79568 152982 79620
rect 152734 79540 152740 79552
rect 152062 79512 152740 79540
rect 152734 79500 152740 79512
rect 152792 79500 152798 79552
rect 143994 79432 144000 79484
rect 144052 79472 144058 79484
rect 151446 79472 151452 79484
rect 144052 79444 151452 79472
rect 144052 79432 144058 79444
rect 151446 79432 151452 79444
rect 151504 79432 151510 79484
rect 153212 79472 153240 79716
rect 153304 79620 153332 79784
rect 153442 79676 153470 79920
rect 153608 79908 153614 79920
rect 153666 79908 153672 79960
rect 153792 79908 153798 79960
rect 153850 79948 153856 79960
rect 153850 79920 153976 79948
rect 153850 79908 153856 79920
rect 153700 79840 153706 79892
rect 153758 79880 153764 79892
rect 153758 79852 153838 79880
rect 153758 79840 153764 79852
rect 153516 79772 153522 79824
rect 153574 79772 153580 79824
rect 153534 79744 153562 79772
rect 153654 79744 153660 79756
rect 153534 79716 153660 79744
rect 153654 79704 153660 79716
rect 153712 79704 153718 79756
rect 153562 79676 153568 79688
rect 153442 79648 153568 79676
rect 153562 79636 153568 79648
rect 153620 79636 153626 79688
rect 153286 79568 153292 79620
rect 153344 79568 153350 79620
rect 153810 79552 153838 79852
rect 153948 79688 153976 79920
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 154086 79688 154114 79908
rect 154160 79772 154166 79824
rect 154218 79772 154224 79824
rect 154178 79744 154206 79772
rect 154178 79716 154252 79744
rect 153930 79636 153936 79688
rect 153988 79636 153994 79688
rect 154086 79648 154120 79688
rect 154114 79636 154120 79648
rect 154172 79636 154178 79688
rect 154224 79552 154252 79716
rect 153810 79512 153844 79552
rect 153838 79500 153844 79512
rect 153896 79500 153902 79552
rect 154206 79500 154212 79552
rect 154264 79500 154270 79552
rect 154500 79472 154528 80056
rect 158318 79988 158622 80016
rect 158318 79960 158346 79988
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 154988 79908 154994 79960
rect 155046 79908 155052 79960
rect 155172 79908 155178 79960
rect 155230 79908 155236 79960
rect 155264 79908 155270 79960
rect 155322 79908 155328 79960
rect 156000 79908 156006 79960
rect 156058 79908 156064 79960
rect 156276 79908 156282 79960
rect 156334 79948 156340 79960
rect 156460 79948 156466 79960
rect 156334 79908 156368 79948
rect 154638 79688 154666 79908
rect 154712 79840 154718 79892
rect 154770 79840 154776 79892
rect 154574 79636 154580 79688
rect 154632 79648 154666 79688
rect 154632 79636 154638 79648
rect 154730 79620 154758 79840
rect 155006 79824 155034 79908
rect 154942 79772 154948 79824
rect 155000 79784 155034 79824
rect 155000 79772 155006 79784
rect 155190 79688 155218 79908
rect 155282 79880 155310 79908
rect 155448 79880 155454 79892
rect 155282 79852 155356 79880
rect 155328 79688 155356 79852
rect 155420 79840 155454 79880
rect 155506 79840 155512 79892
rect 155816 79840 155822 79892
rect 155874 79840 155880 79892
rect 155908 79840 155914 79892
rect 155966 79840 155972 79892
rect 155420 79688 155448 79840
rect 155190 79648 155224 79688
rect 155218 79636 155224 79648
rect 155276 79636 155282 79688
rect 155310 79636 155316 79688
rect 155368 79636 155374 79688
rect 155402 79636 155408 79688
rect 155460 79636 155466 79688
rect 154730 79580 154764 79620
rect 154758 79568 154764 79580
rect 154816 79568 154822 79620
rect 155834 79540 155862 79840
rect 155926 79676 155954 79840
rect 156018 79824 156046 79908
rect 156184 79840 156190 79892
rect 156242 79880 156248 79892
rect 156242 79840 156276 79880
rect 156000 79772 156006 79824
rect 156058 79772 156064 79824
rect 156138 79676 156144 79688
rect 155926 79648 156144 79676
rect 156138 79636 156144 79648
rect 156196 79636 156202 79688
rect 156248 79620 156276 79840
rect 156230 79568 156236 79620
rect 156288 79568 156294 79620
rect 156340 79552 156368 79908
rect 156432 79908 156466 79948
rect 156518 79908 156524 79960
rect 157196 79908 157202 79960
rect 157254 79948 157260 79960
rect 157254 79908 157288 79948
rect 157748 79908 157754 79960
rect 157806 79908 157812 79960
rect 157840 79908 157846 79960
rect 157898 79908 157904 79960
rect 158024 79908 158030 79960
rect 158082 79948 158088 79960
rect 158208 79948 158214 79960
rect 158082 79908 158116 79948
rect 155834 79512 156276 79540
rect 153212 79444 154528 79472
rect 155126 79432 155132 79484
rect 155184 79472 155190 79484
rect 155770 79472 155776 79484
rect 155184 79444 155776 79472
rect 155184 79432 155190 79444
rect 155770 79432 155776 79444
rect 155828 79432 155834 79484
rect 140498 79404 140504 79416
rect 139274 79376 140504 79404
rect 140498 79364 140504 79376
rect 140556 79364 140562 79416
rect 141326 79364 141332 79416
rect 141384 79364 141390 79416
rect 141418 79364 141424 79416
rect 141476 79364 141482 79416
rect 141878 79364 141884 79416
rect 141936 79376 141970 79416
rect 141936 79364 141942 79376
rect 142062 79364 142068 79416
rect 142120 79404 142126 79416
rect 146938 79404 146944 79416
rect 142120 79376 146944 79404
rect 142120 79364 142126 79376
rect 146938 79364 146944 79376
rect 146996 79364 147002 79416
rect 149698 79364 149704 79416
rect 149756 79404 149762 79416
rect 156248 79404 156276 79512
rect 156322 79500 156328 79552
rect 156380 79500 156386 79552
rect 156432 79484 156460 79908
rect 156552 79880 156558 79892
rect 156524 79840 156558 79880
rect 156610 79840 156616 79892
rect 157012 79840 157018 79892
rect 157070 79880 157076 79892
rect 157070 79852 157196 79880
rect 157070 79840 157076 79852
rect 156524 79756 156552 79840
rect 157168 79824 157196 79852
rect 156828 79812 156834 79824
rect 156616 79784 156834 79812
rect 156616 79756 156644 79784
rect 156828 79772 156834 79784
rect 156886 79772 156892 79824
rect 156920 79772 156926 79824
rect 156978 79772 156984 79824
rect 157150 79772 157156 79824
rect 157208 79772 157214 79824
rect 156506 79704 156512 79756
rect 156564 79704 156570 79756
rect 156598 79704 156604 79756
rect 156656 79704 156662 79756
rect 156938 79688 156966 79772
rect 156874 79636 156880 79688
rect 156932 79648 156966 79688
rect 156932 79636 156938 79648
rect 157058 79568 157064 79620
rect 157116 79608 157122 79620
rect 157260 79608 157288 79908
rect 157380 79880 157386 79892
rect 157352 79840 157386 79880
rect 157438 79840 157444 79892
rect 157656 79840 157662 79892
rect 157714 79840 157720 79892
rect 157352 79620 157380 79840
rect 157674 79620 157702 79840
rect 157766 79744 157794 79908
rect 157858 79812 157886 79908
rect 157858 79784 157932 79812
rect 157766 79716 157840 79744
rect 157116 79580 157288 79608
rect 157116 79568 157122 79580
rect 157334 79568 157340 79620
rect 157392 79568 157398 79620
rect 157674 79580 157708 79620
rect 157702 79568 157708 79580
rect 157760 79568 157766 79620
rect 157518 79500 157524 79552
rect 157576 79540 157582 79552
rect 157812 79540 157840 79716
rect 157904 79620 157932 79784
rect 158088 79620 158116 79908
rect 158180 79908 158214 79948
rect 158266 79908 158272 79960
rect 158300 79908 158306 79960
rect 158358 79908 158364 79960
rect 158484 79908 158490 79960
rect 158542 79908 158548 79960
rect 157886 79568 157892 79620
rect 157944 79568 157950 79620
rect 158070 79568 158076 79620
rect 158128 79568 158134 79620
rect 158180 79552 158208 79908
rect 158502 79756 158530 79908
rect 158438 79704 158444 79756
rect 158496 79716 158530 79756
rect 158496 79704 158502 79716
rect 158594 79688 158622 79988
rect 159054 79960 159082 80056
rect 159146 79988 159358 80016
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 158852 79908 158858 79960
rect 158910 79908 158916 79960
rect 159036 79908 159042 79960
rect 159094 79908 159100 79960
rect 158530 79636 158536 79688
rect 158588 79648 158622 79688
rect 158588 79636 158594 79648
rect 158778 79608 158806 79908
rect 158870 79824 158898 79908
rect 158852 79772 158858 79824
rect 158910 79772 158916 79824
rect 159146 79688 159174 79988
rect 159330 79960 159358 79988
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 159496 79908 159502 79960
rect 159554 79908 159560 79960
rect 159588 79908 159594 79960
rect 159646 79948 159652 79960
rect 159646 79920 160278 79948
rect 159646 79908 159652 79920
rect 159082 79636 159088 79688
rect 159140 79648 159174 79688
rect 159238 79676 159266 79908
rect 159404 79840 159410 79892
rect 159462 79840 159468 79892
rect 159422 79688 159450 79840
rect 159238 79648 159312 79676
rect 159140 79636 159146 79648
rect 159284 79620 159312 79648
rect 159358 79636 159364 79688
rect 159416 79648 159450 79688
rect 159416 79636 159422 79648
rect 159174 79608 159180 79620
rect 158778 79580 159180 79608
rect 159174 79568 159180 79580
rect 159232 79568 159238 79620
rect 159266 79568 159272 79620
rect 159324 79568 159330 79620
rect 157576 79512 157840 79540
rect 157576 79500 157582 79512
rect 158162 79500 158168 79552
rect 158220 79500 158226 79552
rect 158898 79500 158904 79552
rect 158956 79540 158962 79552
rect 159514 79540 159542 79908
rect 159680 79880 159686 79892
rect 159652 79840 159686 79880
rect 159738 79840 159744 79892
rect 159956 79840 159962 79892
rect 160014 79840 160020 79892
rect 160140 79840 160146 79892
rect 160198 79840 160204 79892
rect 159652 79676 159680 79840
rect 159726 79704 159732 79756
rect 159784 79744 159790 79756
rect 159974 79744 160002 79840
rect 159784 79716 160002 79744
rect 159784 79704 159790 79716
rect 160002 79676 160008 79688
rect 159652 79648 160008 79676
rect 160002 79636 160008 79648
rect 160060 79636 160066 79688
rect 158956 79512 159542 79540
rect 158956 79500 158962 79512
rect 156414 79432 156420 79484
rect 156472 79432 156478 79484
rect 156966 79404 156972 79416
rect 149756 79376 156184 79404
rect 156248 79376 156972 79404
rect 149756 79364 149762 79376
rect 138290 79336 138296 79348
rect 138170 79308 138296 79336
rect 134576 79296 134582 79308
rect 138290 79296 138296 79308
rect 138348 79296 138354 79348
rect 143506 79308 149836 79336
rect 143506 79268 143534 79308
rect 133846 79240 143534 79268
rect 146938 79160 146944 79212
rect 146996 79200 147002 79212
rect 149698 79200 149704 79212
rect 146996 79172 149704 79200
rect 146996 79160 147002 79172
rect 149698 79160 149704 79172
rect 149756 79160 149762 79212
rect 149808 79200 149836 79308
rect 153746 79296 153752 79348
rect 153804 79336 153810 79348
rect 153930 79336 153936 79348
rect 153804 79308 153936 79336
rect 153804 79296 153810 79308
rect 153930 79296 153936 79308
rect 153988 79296 153994 79348
rect 154850 79296 154856 79348
rect 154908 79336 154914 79348
rect 155126 79336 155132 79348
rect 154908 79308 155132 79336
rect 154908 79296 154914 79308
rect 155126 79296 155132 79308
rect 155184 79296 155190 79348
rect 156156 79336 156184 79376
rect 156966 79364 156972 79376
rect 157024 79364 157030 79416
rect 157610 79364 157616 79416
rect 157668 79404 157674 79416
rect 159910 79404 159916 79416
rect 157668 79376 159916 79404
rect 157668 79364 157674 79376
rect 159910 79364 159916 79376
rect 159968 79364 159974 79416
rect 160158 79404 160186 79840
rect 160250 79620 160278 79920
rect 160324 79908 160330 79960
rect 160382 79908 160388 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160692 79908 160698 79960
rect 160750 79908 160756 79960
rect 161060 79908 161066 79960
rect 161118 79908 161124 79960
rect 161152 79908 161158 79960
rect 161210 79908 161216 79960
rect 161244 79908 161250 79960
rect 161302 79908 161308 79960
rect 160342 79812 160370 79908
rect 160434 79880 160462 79908
rect 160434 79852 160508 79880
rect 160480 79824 160508 79852
rect 160600 79840 160606 79892
rect 160658 79840 160664 79892
rect 160342 79784 160416 79812
rect 160388 79756 160416 79784
rect 160462 79772 160468 79824
rect 160520 79772 160526 79824
rect 160370 79704 160376 79756
rect 160428 79704 160434 79756
rect 160618 79744 160646 79840
rect 160480 79716 160646 79744
rect 160250 79580 160284 79620
rect 160278 79568 160284 79580
rect 160336 79568 160342 79620
rect 160480 79608 160508 79716
rect 160554 79636 160560 79688
rect 160612 79676 160618 79688
rect 160710 79676 160738 79908
rect 160968 79880 160974 79892
rect 160612 79648 160738 79676
rect 160848 79852 160974 79880
rect 160612 79636 160618 79648
rect 160646 79608 160652 79620
rect 160480 79580 160652 79608
rect 160646 79568 160652 79580
rect 160704 79568 160710 79620
rect 160848 79552 160876 79852
rect 160968 79840 160974 79852
rect 161026 79840 161032 79892
rect 161078 79812 161106 79908
rect 161032 79784 161106 79812
rect 161032 79756 161060 79784
rect 161170 79756 161198 79908
rect 161014 79704 161020 79756
rect 161072 79704 161078 79756
rect 161106 79704 161112 79756
rect 161164 79716 161198 79756
rect 161164 79704 161170 79716
rect 161262 79688 161290 79908
rect 161198 79636 161204 79688
rect 161256 79648 161290 79688
rect 161256 79636 161262 79648
rect 161354 79620 161382 80056
rect 161446 80016 161474 80192
rect 161446 79988 162026 80016
rect 161796 79948 161802 79960
rect 161768 79908 161802 79948
rect 161854 79908 161860 79960
rect 161888 79908 161894 79960
rect 161946 79908 161952 79960
rect 161612 79840 161618 79892
rect 161670 79840 161676 79892
rect 161428 79772 161434 79824
rect 161486 79772 161492 79824
rect 161446 79688 161474 79772
rect 161630 79756 161658 79840
rect 161566 79704 161572 79756
rect 161624 79716 161658 79756
rect 161624 79704 161630 79716
rect 161768 79688 161796 79908
rect 161906 79880 161934 79908
rect 161860 79852 161934 79880
rect 161860 79756 161888 79852
rect 161998 79824 162026 79988
rect 162072 79908 162078 79960
rect 162130 79908 162136 79960
rect 161934 79772 161940 79824
rect 161992 79784 162026 79824
rect 161992 79772 161998 79784
rect 162090 79756 162118 79908
rect 162256 79840 162262 79892
rect 162314 79840 162320 79892
rect 162348 79840 162354 79892
rect 162406 79840 162412 79892
rect 162440 79840 162446 79892
rect 162498 79880 162504 79892
rect 162900 79880 162906 79892
rect 162498 79852 162716 79880
rect 162498 79840 162504 79852
rect 161842 79704 161848 79756
rect 161900 79704 161906 79756
rect 162026 79704 162032 79756
rect 162084 79716 162118 79756
rect 162084 79704 162090 79716
rect 162274 79688 162302 79840
rect 162366 79744 162394 79840
rect 162366 79716 162440 79744
rect 161446 79648 161480 79688
rect 161474 79636 161480 79648
rect 161532 79636 161538 79688
rect 161750 79636 161756 79688
rect 161808 79636 161814 79688
rect 162274 79648 162308 79688
rect 162302 79636 162308 79648
rect 162360 79636 162366 79688
rect 161290 79568 161296 79620
rect 161348 79580 161382 79620
rect 161348 79568 161354 79580
rect 162118 79568 162124 79620
rect 162176 79608 162182 79620
rect 162412 79608 162440 79716
rect 162688 79688 162716 79852
rect 162780 79852 162906 79880
rect 162780 79688 162808 79852
rect 162900 79840 162906 79852
rect 162958 79840 162964 79892
rect 163056 79812 163084 80260
rect 163268 79840 163274 79892
rect 163326 79880 163332 79892
rect 163326 79840 163360 79880
rect 163056 79784 163268 79812
rect 163240 79756 163268 79784
rect 163222 79704 163228 79756
rect 163280 79704 163286 79756
rect 163332 79688 163360 79840
rect 163424 79688 163452 80328
rect 174446 80316 174452 80368
rect 174504 80356 174510 80368
rect 180150 80356 180156 80368
rect 174504 80328 180156 80356
rect 174504 80316 174510 80328
rect 180150 80316 180156 80328
rect 180208 80316 180214 80368
rect 164022 80260 171042 80288
rect 164022 80016 164050 80260
rect 163516 79988 164050 80016
rect 167978 79988 168190 80016
rect 162670 79636 162676 79688
rect 162728 79636 162734 79688
rect 162762 79636 162768 79688
rect 162820 79636 162826 79688
rect 163314 79636 163320 79688
rect 163372 79636 163378 79688
rect 163406 79636 163412 79688
rect 163464 79636 163470 79688
rect 162176 79580 162440 79608
rect 162176 79568 162182 79580
rect 162486 79568 162492 79620
rect 162544 79608 162550 79620
rect 163516 79608 163544 79988
rect 163912 79908 163918 79960
rect 163970 79908 163976 79960
rect 164188 79908 164194 79960
rect 164246 79908 164252 79960
rect 164832 79908 164838 79960
rect 164890 79908 164896 79960
rect 164924 79908 164930 79960
rect 164982 79948 164988 79960
rect 164982 79920 165246 79948
rect 164982 79908 164988 79920
rect 163636 79880 163642 79892
rect 162544 79580 163544 79608
rect 163608 79840 163642 79880
rect 163694 79840 163700 79892
rect 163728 79840 163734 79892
rect 163786 79880 163792 79892
rect 163786 79840 163820 79880
rect 162544 79568 162550 79580
rect 160830 79500 160836 79552
rect 160888 79500 160894 79552
rect 161658 79500 161664 79552
rect 161716 79540 161722 79552
rect 162394 79540 162400 79552
rect 161716 79512 162400 79540
rect 161716 79500 161722 79512
rect 162394 79500 162400 79512
rect 162452 79500 162458 79552
rect 163130 79500 163136 79552
rect 163188 79540 163194 79552
rect 163406 79540 163412 79552
rect 163188 79512 163412 79540
rect 163188 79500 163194 79512
rect 163406 79500 163412 79512
rect 163464 79500 163470 79552
rect 163608 79540 163636 79840
rect 163792 79756 163820 79840
rect 163930 79824 163958 79908
rect 163930 79784 163964 79824
rect 163958 79772 163964 79784
rect 164016 79772 164022 79824
rect 163774 79704 163780 79756
rect 163832 79704 163838 79756
rect 164206 79688 164234 79908
rect 164142 79636 164148 79688
rect 164200 79648 164234 79688
rect 164200 79636 164206 79648
rect 164850 79620 164878 79908
rect 164694 79608 164700 79620
rect 164344 79580 164700 79608
rect 164344 79552 164372 79580
rect 164694 79568 164700 79580
rect 164752 79568 164758 79620
rect 164850 79580 164884 79620
rect 164878 79568 164884 79580
rect 164936 79568 164942 79620
rect 163958 79540 163964 79552
rect 163608 79512 163964 79540
rect 163958 79500 163964 79512
rect 164016 79500 164022 79552
rect 164326 79500 164332 79552
rect 164384 79500 164390 79552
rect 165218 79540 165246 79920
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 165844 79908 165850 79960
rect 165902 79908 165908 79960
rect 166028 79908 166034 79960
rect 166086 79908 166092 79960
rect 166304 79908 166310 79960
rect 166362 79908 166368 79960
rect 167408 79908 167414 79960
rect 167466 79948 167472 79960
rect 167466 79908 167500 79948
rect 165770 79812 165798 79908
rect 165724 79784 165798 79812
rect 165724 79676 165752 79784
rect 165862 79756 165890 79908
rect 165936 79840 165942 79892
rect 165994 79840 166000 79892
rect 165798 79704 165804 79756
rect 165856 79716 165890 79756
rect 165954 79744 165982 79840
rect 166046 79824 166074 79908
rect 166028 79772 166034 79824
rect 166086 79772 166092 79824
rect 166120 79772 166126 79824
rect 166178 79772 166184 79824
rect 165954 79716 166028 79744
rect 165856 79704 165862 79716
rect 165890 79676 165896 79688
rect 165724 79648 165896 79676
rect 165890 79636 165896 79648
rect 165948 79636 165954 79688
rect 165706 79568 165712 79620
rect 165764 79608 165770 79620
rect 166000 79608 166028 79716
rect 166138 79688 166166 79772
rect 166322 79688 166350 79908
rect 166948 79840 166954 79892
rect 167006 79840 167012 79892
rect 167132 79840 167138 79892
rect 167190 79840 167196 79892
rect 166138 79648 166172 79688
rect 166166 79636 166172 79648
rect 166224 79636 166230 79688
rect 166322 79648 166356 79688
rect 166350 79636 166356 79648
rect 166408 79636 166414 79688
rect 166966 79620 166994 79840
rect 167150 79812 167178 79840
rect 167362 79812 167368 79824
rect 167150 79784 167368 79812
rect 167362 79772 167368 79784
rect 167420 79772 167426 79824
rect 167178 79636 167184 79688
rect 167236 79676 167242 79688
rect 167472 79676 167500 79908
rect 167236 79648 167500 79676
rect 167978 79676 168006 79988
rect 168052 79908 168058 79960
rect 168110 79908 168116 79960
rect 168070 79744 168098 79908
rect 168162 79892 168190 79988
rect 168328 79908 168334 79960
rect 168386 79948 168392 79960
rect 168386 79920 169064 79948
rect 168386 79908 168392 79920
rect 168144 79840 168150 79892
rect 168202 79840 168208 79892
rect 168512 79880 168518 79892
rect 168392 79852 168518 79880
rect 168392 79756 168420 79852
rect 168512 79840 168518 79852
rect 168570 79840 168576 79892
rect 168604 79840 168610 79892
rect 168662 79840 168668 79892
rect 168696 79840 168702 79892
rect 168754 79840 168760 79892
rect 168070 79716 168236 79744
rect 168208 79688 168236 79716
rect 168374 79704 168380 79756
rect 168432 79704 168438 79756
rect 168466 79704 168472 79756
rect 168524 79744 168530 79756
rect 168622 79744 168650 79840
rect 168524 79716 168650 79744
rect 168524 79704 168530 79716
rect 168714 79688 168742 79840
rect 169036 79688 169064 79920
rect 169524 79908 169530 79960
rect 169582 79908 169588 79960
rect 169542 79688 169570 79908
rect 169984 79880 169990 79892
rect 169956 79840 169990 79880
rect 170042 79840 170048 79892
rect 170352 79840 170358 79892
rect 170410 79840 170416 79892
rect 170812 79840 170818 79892
rect 170870 79840 170876 79892
rect 171014 79880 171042 80260
rect 174630 80248 174636 80300
rect 174688 80288 174694 80300
rect 200114 80288 200120 80300
rect 174688 80260 200120 80288
rect 174688 80248 174694 80260
rect 200114 80248 200120 80260
rect 200172 80248 200178 80300
rect 174446 80220 174452 80232
rect 171520 80192 174452 80220
rect 171520 80152 171548 80192
rect 174446 80180 174452 80192
rect 174504 80180 174510 80232
rect 174538 80180 174544 80232
rect 174596 80220 174602 80232
rect 231854 80220 231860 80232
rect 174596 80192 231860 80220
rect 174596 80180 174602 80192
rect 231854 80180 231860 80192
rect 231912 80180 231918 80232
rect 176010 80152 176016 80164
rect 171474 80124 171548 80152
rect 171658 80124 176016 80152
rect 171474 80084 171502 80124
rect 171290 80056 171502 80084
rect 171290 80016 171318 80056
rect 171658 80016 171686 80124
rect 176010 80112 176016 80124
rect 176068 80112 176074 80164
rect 176102 80112 176108 80164
rect 176160 80152 176166 80164
rect 252554 80152 252560 80164
rect 176160 80124 252560 80152
rect 176160 80112 176166 80124
rect 252554 80112 252560 80124
rect 252612 80112 252618 80164
rect 171106 79988 171318 80016
rect 171428 79988 171686 80016
rect 171750 80056 175136 80084
rect 171106 79960 171134 79988
rect 171088 79908 171094 79960
rect 171146 79908 171152 79960
rect 171272 79908 171278 79960
rect 171330 79948 171336 79960
rect 171428 79948 171456 79988
rect 171750 79948 171778 80056
rect 174538 80016 174544 80028
rect 171330 79920 171456 79948
rect 171658 79920 171778 79948
rect 172164 79988 173112 80016
rect 171330 79908 171336 79920
rect 171014 79852 171088 79880
rect 169956 79688 169984 79840
rect 170370 79744 170398 79840
rect 170720 79772 170726 79824
rect 170778 79812 170784 79824
rect 170830 79812 170858 79840
rect 170778 79784 170858 79812
rect 171060 79812 171088 79852
rect 171548 79840 171554 79892
rect 171606 79880 171612 79892
rect 171658 79880 171686 79920
rect 171606 79852 171686 79880
rect 171606 79840 171612 79852
rect 171732 79840 171738 79892
rect 171790 79840 171796 79892
rect 171226 79812 171232 79824
rect 171060 79784 171232 79812
rect 170778 79772 170784 79784
rect 171226 79772 171232 79784
rect 171284 79772 171290 79824
rect 171364 79772 171370 79824
rect 171422 79772 171428 79824
rect 170858 79744 170864 79756
rect 170370 79716 170864 79744
rect 170858 79704 170864 79716
rect 170916 79704 170922 79756
rect 171382 79744 171410 79772
rect 171502 79744 171508 79756
rect 171382 79716 171508 79744
rect 171502 79704 171508 79716
rect 171560 79704 171566 79756
rect 168098 79676 168104 79688
rect 167978 79648 168104 79676
rect 167236 79636 167242 79648
rect 168098 79636 168104 79648
rect 168156 79636 168162 79688
rect 168190 79636 168196 79688
rect 168248 79636 168254 79688
rect 168650 79636 168656 79688
rect 168708 79648 168742 79688
rect 168708 79636 168714 79648
rect 169018 79636 169024 79688
rect 169076 79636 169082 79688
rect 169478 79636 169484 79688
rect 169536 79648 169570 79688
rect 169536 79636 169542 79648
rect 169938 79636 169944 79688
rect 169996 79636 170002 79688
rect 170628 79636 170634 79688
rect 170686 79676 170692 79688
rect 171134 79676 171140 79688
rect 170686 79648 171140 79676
rect 170686 79636 170692 79648
rect 171134 79636 171140 79648
rect 171192 79636 171198 79688
rect 171594 79636 171600 79688
rect 171652 79676 171658 79688
rect 171750 79676 171778 79840
rect 171652 79648 171778 79676
rect 171652 79636 171658 79648
rect 165764 79580 166028 79608
rect 165764 79568 165770 79580
rect 166074 79568 166080 79620
rect 166132 79608 166138 79620
rect 166626 79608 166632 79620
rect 166132 79580 166632 79608
rect 166132 79568 166138 79580
rect 166626 79568 166632 79580
rect 166684 79568 166690 79620
rect 166902 79568 166908 79620
rect 166960 79580 166994 79620
rect 172164 79608 172192 79988
rect 172376 79948 172382 79960
rect 172348 79908 172382 79948
rect 172434 79908 172440 79960
rect 172348 79824 172376 79908
rect 172560 79840 172566 79892
rect 172618 79840 172624 79892
rect 172652 79840 172658 79892
rect 172710 79840 172716 79892
rect 172928 79840 172934 79892
rect 172986 79840 172992 79892
rect 172330 79772 172336 79824
rect 172388 79772 172394 79824
rect 172578 79756 172606 79840
rect 172514 79704 172520 79756
rect 172572 79716 172606 79756
rect 172572 79704 172578 79716
rect 172670 79620 172698 79840
rect 172946 79676 172974 79840
rect 167840 79580 172192 79608
rect 166960 79568 166966 79580
rect 164712 79512 165246 79540
rect 164712 79484 164740 79512
rect 166534 79500 166540 79552
rect 166592 79540 166598 79552
rect 167840 79540 167868 79580
rect 172238 79568 172244 79620
rect 172296 79608 172302 79620
rect 172296 79580 172560 79608
rect 172296 79568 172302 79580
rect 166592 79512 167868 79540
rect 166592 79500 166598 79512
rect 168742 79500 168748 79552
rect 168800 79540 168806 79552
rect 171502 79540 171508 79552
rect 168800 79512 171508 79540
rect 168800 79500 168806 79512
rect 171502 79500 171508 79512
rect 171560 79500 171566 79552
rect 161842 79432 161848 79484
rect 161900 79472 161906 79484
rect 164510 79472 164516 79484
rect 161900 79444 164516 79472
rect 161900 79432 161906 79444
rect 164510 79432 164516 79444
rect 164568 79432 164574 79484
rect 164694 79432 164700 79484
rect 164752 79432 164758 79484
rect 165062 79432 165068 79484
rect 165120 79472 165126 79484
rect 172422 79472 172428 79484
rect 165120 79444 172428 79472
rect 165120 79432 165126 79444
rect 172422 79432 172428 79444
rect 172480 79432 172486 79484
rect 172532 79472 172560 79580
rect 172606 79568 172612 79620
rect 172664 79580 172698 79620
rect 172900 79648 172974 79676
rect 172664 79568 172670 79580
rect 172698 79472 172704 79484
rect 172532 79444 172704 79472
rect 172698 79432 172704 79444
rect 172756 79432 172762 79484
rect 172900 79472 172928 79648
rect 173084 79608 173112 79988
rect 173590 79988 174544 80016
rect 173590 79960 173618 79988
rect 174538 79976 174544 79988
rect 174596 79976 174602 80028
rect 175108 80016 175136 80056
rect 175182 80044 175188 80096
rect 175240 80084 175246 80096
rect 430574 80084 430580 80096
rect 175240 80056 430580 80084
rect 175240 80044 175246 80056
rect 430574 80044 430580 80056
rect 430632 80044 430638 80096
rect 178402 80016 178408 80028
rect 175108 79988 178408 80016
rect 178402 79976 178408 79988
rect 178460 79976 178466 80028
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173940 79908 173946 79960
rect 173998 79908 174004 79960
rect 173204 79840 173210 79892
rect 173262 79880 173268 79892
rect 173262 79840 173296 79880
rect 173268 79756 173296 79840
rect 173682 79824 173710 79908
rect 173664 79772 173670 79824
rect 173722 79772 173728 79824
rect 173250 79704 173256 79756
rect 173308 79704 173314 79756
rect 173958 79744 173986 79908
rect 174124 79840 174130 79892
rect 174182 79840 174188 79892
rect 173636 79716 173986 79744
rect 174142 79756 174170 79840
rect 174142 79716 174176 79756
rect 173636 79688 173664 79716
rect 174170 79704 174176 79716
rect 174228 79704 174234 79756
rect 173618 79636 173624 79688
rect 173676 79636 173682 79688
rect 173802 79608 173808 79620
rect 173084 79580 173808 79608
rect 173802 79568 173808 79580
rect 173860 79568 173866 79620
rect 174722 79472 174728 79484
rect 172900 79444 174728 79472
rect 174722 79432 174728 79444
rect 174780 79432 174786 79484
rect 171778 79404 171784 79416
rect 160158 79376 171784 79404
rect 171778 79364 171784 79376
rect 171836 79364 171842 79416
rect 172146 79364 172152 79416
rect 172204 79404 172210 79416
rect 175274 79404 175280 79416
rect 172204 79376 175280 79404
rect 172204 79364 172210 79376
rect 175274 79364 175280 79376
rect 175332 79364 175338 79416
rect 178034 79404 178040 79416
rect 176626 79376 178040 79404
rect 159634 79336 159640 79348
rect 156156 79308 159640 79336
rect 159634 79296 159640 79308
rect 159692 79296 159698 79348
rect 161934 79296 161940 79348
rect 161992 79336 161998 79348
rect 163406 79336 163412 79348
rect 161992 79308 163412 79336
rect 161992 79296 161998 79308
rect 163406 79296 163412 79308
rect 163464 79296 163470 79348
rect 163792 79308 165200 79336
rect 150342 79228 150348 79280
rect 150400 79268 150406 79280
rect 150400 79240 162808 79268
rect 150400 79228 150406 79240
rect 162780 79200 162808 79240
rect 163792 79200 163820 79308
rect 164510 79228 164516 79280
rect 164568 79268 164574 79280
rect 165062 79268 165068 79280
rect 164568 79240 165068 79268
rect 164568 79228 164574 79240
rect 165062 79228 165068 79240
rect 165120 79228 165126 79280
rect 165172 79268 165200 79308
rect 166626 79296 166632 79348
rect 166684 79336 166690 79348
rect 166994 79336 167000 79348
rect 166684 79308 167000 79336
rect 166684 79296 166690 79308
rect 166994 79296 167000 79308
rect 167052 79296 167058 79348
rect 167454 79296 167460 79348
rect 167512 79336 167518 79348
rect 176626 79336 176654 79376
rect 178034 79364 178040 79376
rect 178092 79364 178098 79416
rect 167512 79308 176654 79336
rect 167512 79296 167518 79308
rect 179414 79296 179420 79348
rect 179472 79336 179478 79348
rect 580442 79336 580448 79348
rect 179472 79308 580448 79336
rect 179472 79296 179478 79308
rect 580442 79296 580448 79308
rect 580500 79296 580506 79348
rect 174170 79268 174176 79280
rect 165172 79240 174176 79268
rect 174170 79228 174176 79240
rect 174228 79228 174234 79280
rect 174262 79200 174268 79212
rect 149808 79172 162440 79200
rect 162780 79172 163820 79200
rect 164206 79172 174268 79200
rect 120442 79092 120448 79144
rect 120500 79132 120506 79144
rect 150342 79132 150348 79144
rect 120500 79104 138704 79132
rect 120500 79092 120506 79104
rect 118666 79036 133874 79064
rect 5074 78820 5080 78872
rect 5132 78860 5138 78872
rect 118666 78860 118694 79036
rect 133846 78928 133874 79036
rect 138676 78996 138704 79104
rect 138860 79104 150348 79132
rect 138860 78996 138888 79104
rect 150342 79092 150348 79104
rect 150400 79092 150406 79144
rect 151446 79092 151452 79144
rect 151504 79132 151510 79144
rect 161842 79132 161848 79144
rect 151504 79104 161848 79132
rect 151504 79092 151510 79104
rect 161842 79092 161848 79104
rect 161900 79092 161906 79144
rect 145190 79024 145196 79076
rect 145248 79064 145254 79076
rect 147582 79064 147588 79076
rect 145248 79036 147588 79064
rect 145248 79024 145254 79036
rect 147582 79024 147588 79036
rect 147640 79024 147646 79076
rect 148962 79024 148968 79076
rect 149020 79064 149026 79076
rect 149020 79036 159404 79064
rect 149020 79024 149026 79036
rect 157242 78996 157248 79008
rect 138676 78968 138888 78996
rect 143506 78968 157248 78996
rect 143506 78928 143534 78968
rect 157242 78956 157248 78968
rect 157300 78956 157306 79008
rect 159376 78996 159404 79036
rect 160554 79024 160560 79076
rect 160612 79064 160618 79076
rect 161290 79064 161296 79076
rect 160612 79036 161296 79064
rect 160612 79024 160618 79036
rect 161290 79024 161296 79036
rect 161348 79024 161354 79076
rect 162412 79064 162440 79172
rect 163498 79092 163504 79144
rect 163556 79132 163562 79144
rect 164206 79132 164234 79172
rect 174262 79160 174268 79172
rect 174320 79160 174326 79212
rect 166534 79132 166540 79144
rect 163556 79104 164234 79132
rect 164988 79104 166540 79132
rect 163556 79092 163562 79104
rect 164988 79064 165016 79104
rect 166534 79092 166540 79104
rect 166592 79092 166598 79144
rect 166902 79092 166908 79144
rect 166960 79132 166966 79144
rect 195974 79132 195980 79144
rect 166960 79104 195980 79132
rect 166960 79092 166966 79104
rect 195974 79092 195980 79104
rect 196032 79092 196038 79144
rect 162412 79036 165016 79064
rect 165062 79024 165068 79076
rect 165120 79064 165126 79076
rect 249794 79064 249800 79076
rect 165120 79036 249800 79064
rect 165120 79024 165126 79036
rect 249794 79024 249800 79036
rect 249852 79024 249858 79076
rect 164510 78996 164516 79008
rect 159376 78968 164516 78996
rect 164510 78956 164516 78968
rect 164568 78956 164574 79008
rect 165614 78956 165620 79008
rect 165672 78996 165678 79008
rect 165672 78968 166488 78996
rect 165672 78956 165678 78968
rect 133846 78900 143534 78928
rect 144454 78888 144460 78940
rect 144512 78928 144518 78940
rect 146938 78928 146944 78940
rect 144512 78900 146944 78928
rect 144512 78888 144518 78900
rect 146938 78888 146944 78900
rect 146996 78888 147002 78940
rect 155034 78888 155040 78940
rect 155092 78928 155098 78940
rect 155494 78928 155500 78940
rect 155092 78900 155500 78928
rect 155092 78888 155098 78900
rect 155494 78888 155500 78900
rect 155552 78888 155558 78940
rect 157702 78888 157708 78940
rect 157760 78928 157766 78940
rect 157978 78928 157984 78940
rect 157760 78900 157984 78928
rect 157760 78888 157766 78900
rect 157978 78888 157984 78900
rect 158036 78888 158042 78940
rect 159358 78888 159364 78940
rect 159416 78928 159422 78940
rect 160278 78928 160284 78940
rect 159416 78900 160284 78928
rect 159416 78888 159422 78900
rect 160278 78888 160284 78900
rect 160336 78888 160342 78940
rect 161658 78888 161664 78940
rect 161716 78928 161722 78940
rect 162210 78928 162216 78940
rect 161716 78900 162216 78928
rect 161716 78888 161722 78900
rect 162210 78888 162216 78900
rect 162268 78888 162274 78940
rect 162578 78888 162584 78940
rect 162636 78928 162642 78940
rect 162946 78928 162952 78940
rect 162636 78900 162952 78928
rect 162636 78888 162642 78900
rect 162946 78888 162952 78900
rect 163004 78888 163010 78940
rect 164234 78888 164240 78940
rect 164292 78928 164298 78940
rect 164786 78928 164792 78940
rect 164292 78900 164792 78928
rect 164292 78888 164298 78900
rect 164786 78888 164792 78900
rect 164844 78888 164850 78940
rect 165706 78888 165712 78940
rect 165764 78928 165770 78940
rect 166074 78928 166080 78940
rect 165764 78900 166080 78928
rect 165764 78888 165770 78900
rect 166074 78888 166080 78900
rect 166132 78888 166138 78940
rect 166460 78928 166488 78968
rect 166534 78956 166540 79008
rect 166592 78996 166598 79008
rect 166592 78968 166948 78996
rect 166592 78956 166598 78968
rect 166920 78928 166948 78968
rect 166994 78956 167000 79008
rect 167052 78996 167058 79008
rect 171318 78996 171324 79008
rect 167052 78968 171324 78996
rect 167052 78956 167058 78968
rect 171318 78956 171324 78968
rect 171376 78956 171382 79008
rect 171686 78956 171692 79008
rect 171744 78996 171750 79008
rect 213914 78996 213920 79008
rect 171744 78968 213920 78996
rect 171744 78956 171750 78968
rect 213914 78956 213920 78968
rect 213972 78956 213978 79008
rect 267734 78928 267740 78940
rect 166460 78900 166856 78928
rect 166920 78900 267740 78928
rect 5132 78832 118694 78860
rect 5132 78820 5138 78832
rect 134058 78820 134064 78872
rect 134116 78860 134122 78872
rect 143994 78860 144000 78872
rect 134116 78832 144000 78860
rect 134116 78820 134122 78832
rect 143994 78820 144000 78832
rect 144052 78820 144058 78872
rect 145190 78820 145196 78872
rect 145248 78860 145254 78872
rect 145650 78860 145656 78872
rect 145248 78832 145656 78860
rect 145248 78820 145254 78832
rect 145650 78820 145656 78832
rect 145708 78820 145714 78872
rect 148318 78820 148324 78872
rect 148376 78860 148382 78872
rect 148502 78860 148508 78872
rect 148376 78832 148508 78860
rect 148376 78820 148382 78832
rect 148502 78820 148508 78832
rect 148560 78820 148566 78872
rect 159174 78820 159180 78872
rect 159232 78860 159238 78872
rect 166626 78860 166632 78872
rect 159232 78832 166632 78860
rect 159232 78820 159238 78832
rect 166626 78820 166632 78832
rect 166684 78820 166690 78872
rect 157610 78752 157616 78804
rect 157668 78792 157674 78804
rect 158070 78792 158076 78804
rect 157668 78764 158076 78792
rect 157668 78752 157674 78764
rect 158070 78752 158076 78764
rect 158128 78752 158134 78804
rect 160186 78752 160192 78804
rect 160244 78792 160250 78804
rect 160922 78792 160928 78804
rect 160244 78764 160928 78792
rect 160244 78752 160250 78764
rect 160922 78752 160928 78764
rect 160980 78752 160986 78804
rect 161566 78752 161572 78804
rect 161624 78792 161630 78804
rect 161934 78792 161940 78804
rect 161624 78764 161940 78792
rect 161624 78752 161630 78764
rect 161934 78752 161940 78764
rect 161992 78752 161998 78804
rect 162210 78752 162216 78804
rect 162268 78792 162274 78804
rect 165062 78792 165068 78804
rect 162268 78764 165068 78792
rect 162268 78752 162274 78764
rect 165062 78752 165068 78764
rect 165120 78752 165126 78804
rect 165798 78752 165804 78804
rect 165856 78792 165862 78804
rect 166074 78792 166080 78804
rect 165856 78764 166080 78792
rect 165856 78752 165862 78764
rect 166074 78752 166080 78764
rect 166132 78752 166138 78804
rect 166828 78792 166856 78900
rect 267734 78888 267740 78900
rect 267792 78888 267798 78940
rect 166994 78820 167000 78872
rect 167052 78860 167058 78872
rect 171870 78860 171876 78872
rect 167052 78832 171876 78860
rect 167052 78820 167058 78832
rect 171870 78820 171876 78832
rect 171928 78820 171934 78872
rect 172514 78820 172520 78872
rect 172572 78860 172578 78872
rect 293218 78860 293224 78872
rect 172572 78832 293224 78860
rect 172572 78820 172578 78832
rect 293218 78820 293224 78832
rect 293276 78820 293282 78872
rect 168282 78792 168288 78804
rect 166828 78764 168288 78792
rect 168282 78752 168288 78764
rect 168340 78752 168346 78804
rect 170490 78752 170496 78804
rect 170548 78792 170554 78804
rect 170858 78792 170864 78804
rect 170548 78764 170864 78792
rect 170548 78752 170554 78764
rect 170858 78752 170864 78764
rect 170916 78752 170922 78804
rect 171778 78752 171784 78804
rect 171836 78792 171842 78804
rect 444374 78792 444380 78804
rect 171836 78764 444380 78792
rect 171836 78752 171842 78764
rect 444374 78752 444380 78764
rect 444432 78752 444438 78804
rect 115290 78684 115296 78736
rect 115348 78724 115354 78736
rect 115348 78696 115980 78724
rect 115348 78684 115354 78696
rect 115952 78656 115980 78696
rect 131574 78684 131580 78736
rect 131632 78724 131638 78736
rect 133874 78724 133880 78736
rect 131632 78696 133880 78724
rect 131632 78684 131638 78696
rect 133874 78684 133880 78696
rect 133932 78684 133938 78736
rect 146846 78684 146852 78736
rect 146904 78724 146910 78736
rect 147306 78724 147312 78736
rect 146904 78696 147312 78724
rect 146904 78684 146910 78696
rect 147306 78684 147312 78696
rect 147364 78684 147370 78736
rect 147950 78684 147956 78736
rect 148008 78724 148014 78736
rect 148134 78724 148140 78736
rect 148008 78696 148140 78724
rect 148008 78684 148014 78696
rect 148134 78684 148140 78696
rect 148192 78684 148198 78736
rect 148318 78684 148324 78736
rect 148376 78724 148382 78736
rect 148686 78724 148692 78736
rect 148376 78696 148692 78724
rect 148376 78684 148382 78696
rect 148686 78684 148692 78696
rect 148744 78684 148750 78736
rect 159174 78724 159180 78736
rect 154546 78696 159180 78724
rect 119982 78656 119988 78668
rect 115952 78628 119988 78656
rect 119982 78616 119988 78628
rect 120040 78616 120046 78668
rect 145650 78616 145656 78668
rect 145708 78656 145714 78668
rect 146018 78656 146024 78668
rect 145708 78628 146024 78656
rect 145708 78616 145714 78628
rect 146018 78616 146024 78628
rect 146076 78616 146082 78668
rect 146386 78616 146392 78668
rect 146444 78656 146450 78668
rect 146754 78656 146760 78668
rect 146444 78628 146760 78656
rect 146444 78616 146450 78628
rect 146754 78616 146760 78628
rect 146812 78616 146818 78668
rect 147582 78616 147588 78668
rect 147640 78656 147646 78668
rect 154546 78656 154574 78696
rect 159174 78684 159180 78696
rect 159232 78684 159238 78736
rect 161842 78684 161848 78736
rect 161900 78724 161906 78736
rect 162118 78724 162124 78736
rect 161900 78696 162124 78724
rect 161900 78684 161906 78696
rect 162118 78684 162124 78696
rect 162176 78684 162182 78736
rect 164510 78684 164516 78736
rect 164568 78724 164574 78736
rect 166534 78724 166540 78736
rect 164568 78696 166540 78724
rect 164568 78684 164574 78696
rect 166534 78684 166540 78696
rect 166592 78684 166598 78736
rect 168650 78684 168656 78736
rect 168708 78724 168714 78736
rect 554774 78724 554780 78736
rect 168708 78696 554780 78724
rect 168708 78684 168714 78696
rect 554774 78684 554780 78696
rect 554832 78684 554838 78736
rect 147640 78628 154574 78656
rect 147640 78616 147646 78628
rect 157886 78616 157892 78668
rect 157944 78656 157950 78668
rect 158070 78656 158076 78668
rect 157944 78628 158076 78656
rect 157944 78616 157950 78628
rect 158070 78616 158076 78628
rect 158128 78616 158134 78668
rect 160554 78616 160560 78668
rect 160612 78656 160618 78668
rect 160830 78656 160836 78668
rect 160612 78628 160836 78656
rect 160612 78616 160618 78628
rect 160830 78616 160836 78628
rect 160888 78616 160894 78668
rect 160922 78616 160928 78668
rect 160980 78656 160986 78668
rect 170858 78656 170864 78668
rect 160980 78628 170864 78656
rect 160980 78616 160986 78628
rect 170858 78616 170864 78628
rect 170916 78616 170922 78668
rect 171778 78656 171784 78668
rect 171336 78628 171784 78656
rect 139670 78548 139676 78600
rect 139728 78588 139734 78600
rect 171336 78588 171364 78628
rect 171778 78616 171784 78628
rect 171836 78616 171842 78668
rect 171962 78616 171968 78668
rect 172020 78656 172026 78668
rect 179414 78656 179420 78668
rect 172020 78628 179420 78656
rect 172020 78616 172026 78628
rect 179414 78616 179420 78628
rect 179472 78616 179478 78668
rect 139728 78560 171364 78588
rect 139728 78548 139734 78560
rect 172422 78548 172428 78600
rect 172480 78588 172486 78600
rect 173618 78588 173624 78600
rect 172480 78560 173624 78588
rect 172480 78548 172486 78560
rect 173618 78548 173624 78560
rect 173676 78548 173682 78600
rect 178954 78588 178960 78600
rect 173866 78560 178960 78588
rect 128630 78480 128636 78532
rect 128688 78520 128694 78532
rect 131206 78520 131212 78532
rect 128688 78492 131212 78520
rect 128688 78480 128694 78492
rect 131206 78480 131212 78492
rect 131264 78480 131270 78532
rect 140774 78480 140780 78532
rect 140832 78520 140838 78532
rect 166902 78520 166908 78532
rect 140832 78492 166908 78520
rect 140832 78480 140838 78492
rect 166902 78480 166908 78492
rect 166960 78480 166966 78532
rect 171686 78520 171692 78532
rect 170784 78492 171692 78520
rect 142614 78412 142620 78464
rect 142672 78452 142678 78464
rect 160922 78452 160928 78464
rect 142672 78424 160928 78452
rect 142672 78412 142678 78424
rect 160922 78412 160928 78424
rect 160980 78412 160986 78464
rect 161198 78412 161204 78464
rect 161256 78452 161262 78464
rect 163130 78452 163136 78464
rect 161256 78424 163136 78452
rect 161256 78412 161262 78424
rect 163130 78412 163136 78424
rect 163188 78412 163194 78464
rect 170784 78452 170812 78492
rect 171686 78480 171692 78492
rect 171744 78480 171750 78532
rect 172054 78480 172060 78532
rect 172112 78520 172118 78532
rect 173866 78520 173894 78560
rect 178954 78548 178960 78560
rect 179012 78548 179018 78600
rect 172112 78492 173894 78520
rect 172112 78480 172118 78492
rect 163700 78424 163958 78452
rect 125318 78344 125324 78396
rect 125376 78384 125382 78396
rect 125594 78384 125600 78396
rect 125376 78356 125600 78384
rect 125376 78344 125382 78356
rect 125594 78344 125600 78356
rect 125652 78344 125658 78396
rect 142246 78344 142252 78396
rect 142304 78384 142310 78396
rect 163700 78384 163728 78424
rect 142304 78356 163728 78384
rect 163930 78384 163958 78424
rect 164206 78424 170812 78452
rect 164206 78384 164234 78424
rect 171226 78412 171232 78464
rect 171284 78452 171290 78464
rect 175182 78452 175188 78464
rect 171284 78424 175188 78452
rect 171284 78412 171290 78424
rect 175182 78412 175188 78424
rect 175240 78412 175246 78464
rect 163930 78356 164234 78384
rect 142304 78344 142310 78356
rect 164786 78344 164792 78396
rect 164844 78384 164850 78396
rect 166994 78384 167000 78396
rect 164844 78356 167000 78384
rect 164844 78344 164850 78356
rect 166994 78344 167000 78356
rect 167052 78344 167058 78396
rect 167086 78344 167092 78396
rect 167144 78384 167150 78396
rect 173158 78384 173164 78396
rect 167144 78356 173164 78384
rect 167144 78344 167150 78356
rect 173158 78344 173164 78356
rect 173216 78344 173222 78396
rect 120810 78276 120816 78328
rect 120868 78316 120874 78328
rect 129090 78316 129096 78328
rect 120868 78288 129096 78316
rect 120868 78276 120874 78288
rect 129090 78276 129096 78288
rect 129148 78276 129154 78328
rect 131206 78276 131212 78328
rect 131264 78316 131270 78328
rect 131942 78316 131948 78328
rect 131264 78288 131948 78316
rect 131264 78276 131270 78288
rect 131942 78276 131948 78288
rect 132000 78276 132006 78328
rect 152642 78276 152648 78328
rect 152700 78316 152706 78328
rect 160922 78316 160928 78328
rect 152700 78288 160928 78316
rect 152700 78276 152706 78288
rect 160922 78276 160928 78288
rect 160980 78276 160986 78328
rect 161106 78276 161112 78328
rect 161164 78316 161170 78328
rect 247678 78316 247684 78328
rect 161164 78288 247684 78316
rect 161164 78276 161170 78288
rect 247678 78276 247684 78288
rect 247736 78276 247742 78328
rect 125226 78208 125232 78260
rect 125284 78248 125290 78260
rect 132954 78248 132960 78260
rect 125284 78220 132960 78248
rect 125284 78208 125290 78220
rect 132954 78208 132960 78220
rect 133012 78208 133018 78260
rect 154206 78208 154212 78260
rect 154264 78248 154270 78260
rect 154666 78248 154672 78260
rect 154264 78220 154672 78248
rect 154264 78208 154270 78220
rect 154666 78208 154672 78220
rect 154724 78208 154730 78260
rect 160738 78208 160744 78260
rect 160796 78248 160802 78260
rect 161290 78248 161296 78260
rect 160796 78220 161296 78248
rect 160796 78208 160802 78220
rect 161290 78208 161296 78220
rect 161348 78208 161354 78260
rect 162394 78208 162400 78260
rect 162452 78248 162458 78260
rect 253198 78248 253204 78260
rect 162452 78220 253204 78248
rect 162452 78208 162458 78220
rect 253198 78208 253204 78220
rect 253256 78208 253262 78260
rect 89714 78140 89720 78192
rect 89772 78180 89778 78192
rect 132402 78180 132408 78192
rect 89772 78152 132408 78180
rect 89772 78140 89778 78152
rect 132402 78140 132408 78152
rect 132460 78140 132466 78192
rect 133966 78140 133972 78192
rect 134024 78180 134030 78192
rect 134426 78180 134432 78192
rect 134024 78152 134432 78180
rect 134024 78140 134030 78152
rect 134426 78140 134432 78152
rect 134484 78140 134490 78192
rect 155126 78140 155132 78192
rect 155184 78180 155190 78192
rect 161014 78180 161020 78192
rect 155184 78152 161020 78180
rect 155184 78140 155190 78152
rect 161014 78140 161020 78152
rect 161072 78140 161078 78192
rect 162946 78140 162952 78192
rect 163004 78180 163010 78192
rect 163590 78180 163596 78192
rect 163004 78152 163596 78180
rect 163004 78140 163010 78152
rect 163590 78140 163596 78152
rect 163648 78140 163654 78192
rect 165338 78140 165344 78192
rect 165396 78180 165402 78192
rect 168742 78180 168748 78192
rect 165396 78152 168748 78180
rect 165396 78140 165402 78152
rect 168742 78140 168748 78152
rect 168800 78140 168806 78192
rect 170122 78140 170128 78192
rect 170180 78180 170186 78192
rect 170674 78180 170680 78192
rect 170180 78152 170680 78180
rect 170180 78140 170186 78152
rect 170674 78140 170680 78152
rect 170732 78140 170738 78192
rect 171042 78140 171048 78192
rect 171100 78180 171106 78192
rect 322198 78180 322204 78192
rect 171100 78152 322204 78180
rect 171100 78140 171106 78152
rect 322198 78140 322204 78152
rect 322256 78140 322262 78192
rect 57238 78072 57244 78124
rect 57296 78112 57302 78124
rect 126974 78112 126980 78124
rect 57296 78084 126980 78112
rect 57296 78072 57302 78084
rect 126974 78072 126980 78084
rect 127032 78072 127038 78124
rect 140866 78072 140872 78124
rect 140924 78112 140930 78124
rect 140924 78084 150296 78112
rect 140924 78072 140930 78084
rect 150268 78056 150296 78084
rect 159634 78072 159640 78124
rect 159692 78112 159698 78124
rect 162118 78112 162124 78124
rect 159692 78084 162124 78112
rect 159692 78072 159698 78084
rect 162118 78072 162124 78084
rect 162176 78072 162182 78124
rect 162302 78072 162308 78124
rect 162360 78112 162366 78124
rect 471974 78112 471980 78124
rect 162360 78084 471980 78112
rect 162360 78072 162366 78084
rect 471974 78072 471980 78084
rect 472032 78072 472038 78124
rect 46198 78004 46204 78056
rect 46256 78044 46262 78056
rect 126330 78044 126336 78056
rect 46256 78016 126336 78044
rect 46256 78004 46262 78016
rect 126330 78004 126336 78016
rect 126388 78004 126394 78056
rect 129090 78004 129096 78056
rect 129148 78044 129154 78056
rect 129458 78044 129464 78056
rect 129148 78016 129464 78044
rect 129148 78004 129154 78016
rect 129458 78004 129464 78016
rect 129516 78004 129522 78056
rect 129642 78004 129648 78056
rect 129700 78044 129706 78056
rect 129826 78044 129832 78056
rect 129700 78016 129832 78044
rect 129700 78004 129706 78016
rect 129826 78004 129832 78016
rect 129884 78004 129890 78056
rect 134426 78004 134432 78056
rect 134484 78044 134490 78056
rect 135162 78044 135168 78056
rect 134484 78016 135168 78044
rect 134484 78004 134490 78016
rect 135162 78004 135168 78016
rect 135220 78004 135226 78056
rect 140314 78004 140320 78056
rect 140372 78044 140378 78056
rect 148686 78044 148692 78056
rect 140372 78016 148692 78044
rect 140372 78004 140378 78016
rect 148686 78004 148692 78016
rect 148744 78004 148750 78056
rect 150250 78004 150256 78056
rect 150308 78004 150314 78056
rect 154298 78004 154304 78056
rect 154356 78044 154362 78056
rect 162394 78044 162400 78056
rect 154356 78016 162400 78044
rect 154356 78004 154362 78016
rect 162394 78004 162400 78016
rect 162452 78004 162458 78056
rect 162762 78004 162768 78056
rect 162820 78044 162826 78056
rect 480254 78044 480260 78056
rect 162820 78016 480260 78044
rect 162820 78004 162826 78016
rect 480254 78004 480260 78016
rect 480312 78004 480318 78056
rect 22738 77936 22744 77988
rect 22796 77976 22802 77988
rect 122926 77976 122932 77988
rect 22796 77948 122932 77976
rect 22796 77936 22802 77948
rect 122926 77936 122932 77948
rect 122984 77936 122990 77988
rect 125134 77936 125140 77988
rect 125192 77976 125198 77988
rect 127066 77976 127072 77988
rect 125192 77948 127072 77976
rect 125192 77936 125198 77948
rect 127066 77936 127072 77948
rect 127124 77936 127130 77988
rect 128998 77936 129004 77988
rect 129056 77976 129062 77988
rect 131390 77976 131396 77988
rect 129056 77948 131396 77976
rect 129056 77936 129062 77948
rect 131390 77936 131396 77948
rect 131448 77936 131454 77988
rect 132218 77936 132224 77988
rect 132276 77976 132282 77988
rect 132678 77976 132684 77988
rect 132276 77948 132684 77976
rect 132276 77936 132282 77948
rect 132678 77936 132684 77948
rect 132736 77936 132742 77988
rect 133874 77936 133880 77988
rect 133932 77976 133938 77988
rect 135898 77976 135904 77988
rect 133932 77948 135904 77976
rect 133932 77936 133938 77948
rect 135898 77936 135904 77948
rect 135956 77936 135962 77988
rect 156138 77936 156144 77988
rect 156196 77976 156202 77988
rect 156196 77948 158714 77976
rect 156196 77936 156202 77948
rect 125318 77868 125324 77920
rect 125376 77908 125382 77920
rect 133414 77908 133420 77920
rect 125376 77880 133420 77908
rect 125376 77868 125382 77880
rect 133414 77868 133420 77880
rect 133472 77868 133478 77920
rect 135438 77868 135444 77920
rect 135496 77908 135502 77920
rect 136542 77908 136548 77920
rect 135496 77880 136548 77908
rect 135496 77868 135502 77880
rect 136542 77868 136548 77880
rect 136600 77868 136606 77920
rect 158686 77908 158714 77948
rect 160646 77936 160652 77988
rect 160704 77976 160710 77988
rect 160704 77948 166994 77976
rect 160704 77936 160710 77948
rect 162302 77908 162308 77920
rect 158686 77880 162308 77908
rect 162302 77868 162308 77880
rect 162360 77868 162366 77920
rect 163222 77868 163228 77920
rect 163280 77908 163286 77920
rect 164050 77908 164056 77920
rect 163280 77880 164056 77908
rect 163280 77868 163286 77880
rect 164050 77868 164056 77880
rect 164108 77868 164114 77920
rect 164786 77868 164792 77920
rect 164844 77908 164850 77920
rect 165154 77908 165160 77920
rect 164844 77880 165160 77908
rect 164844 77868 164850 77880
rect 165154 77868 165160 77880
rect 165212 77868 165218 77920
rect 166966 77908 166994 77948
rect 168742 77936 168748 77988
rect 168800 77976 168806 77988
rect 498194 77976 498200 77988
rect 168800 77948 498200 77976
rect 168800 77936 168806 77948
rect 498194 77936 498200 77948
rect 498252 77936 498258 77988
rect 180058 77908 180064 77920
rect 166966 77880 180064 77908
rect 180058 77868 180064 77880
rect 180116 77868 180122 77920
rect 126974 77800 126980 77852
rect 127032 77840 127038 77852
rect 129366 77840 129372 77852
rect 127032 77812 129372 77840
rect 127032 77800 127038 77812
rect 129366 77800 129372 77812
rect 129424 77800 129430 77852
rect 129734 77800 129740 77852
rect 129792 77840 129798 77852
rect 130562 77840 130568 77852
rect 129792 77812 130568 77840
rect 129792 77800 129798 77812
rect 130562 77800 130568 77812
rect 130620 77800 130626 77852
rect 133046 77800 133052 77852
rect 133104 77840 133110 77852
rect 133230 77840 133236 77852
rect 133104 77812 133236 77840
rect 133104 77800 133110 77812
rect 133230 77800 133236 77812
rect 133288 77800 133294 77852
rect 151538 77800 151544 77852
rect 151596 77840 151602 77852
rect 156138 77840 156144 77852
rect 151596 77812 156144 77840
rect 151596 77800 151602 77812
rect 156138 77800 156144 77812
rect 156196 77800 156202 77852
rect 158622 77800 158628 77852
rect 158680 77840 158686 77852
rect 174538 77840 174544 77852
rect 158680 77812 174544 77840
rect 158680 77800 158686 77812
rect 174538 77800 174544 77812
rect 174596 77800 174602 77852
rect 123478 77732 123484 77784
rect 123536 77772 123542 77784
rect 134886 77772 134892 77784
rect 123536 77744 134892 77772
rect 123536 77732 123542 77744
rect 134886 77732 134892 77744
rect 134944 77732 134950 77784
rect 159266 77732 159272 77784
rect 159324 77772 159330 77784
rect 175918 77772 175924 77784
rect 159324 77744 175924 77772
rect 159324 77732 159330 77744
rect 175918 77732 175924 77744
rect 175976 77732 175982 77784
rect 122558 77664 122564 77716
rect 122616 77704 122622 77716
rect 127618 77704 127624 77716
rect 122616 77676 127624 77704
rect 122616 77664 122622 77676
rect 127618 77664 127624 77676
rect 127676 77664 127682 77716
rect 132770 77664 132776 77716
rect 132828 77704 132834 77716
rect 133230 77704 133236 77716
rect 132828 77676 133236 77704
rect 132828 77664 132834 77676
rect 133230 77664 133236 77676
rect 133288 77664 133294 77716
rect 138014 77664 138020 77716
rect 138072 77704 138078 77716
rect 139026 77704 139032 77716
rect 138072 77676 139032 77704
rect 138072 77664 138078 77676
rect 139026 77664 139032 77676
rect 139084 77664 139090 77716
rect 139302 77664 139308 77716
rect 139360 77704 139366 77716
rect 139360 77676 154712 77704
rect 139360 77664 139366 77676
rect 129366 77596 129372 77648
rect 129424 77636 129430 77648
rect 130194 77636 130200 77648
rect 129424 77608 130200 77636
rect 129424 77596 129430 77608
rect 130194 77596 130200 77608
rect 130252 77596 130258 77648
rect 143626 77596 143632 77648
rect 143684 77636 143690 77648
rect 153286 77636 153292 77648
rect 143684 77608 153292 77636
rect 143684 77596 143690 77608
rect 153286 77596 153292 77608
rect 153344 77596 153350 77648
rect 131666 77528 131672 77580
rect 131724 77568 131730 77580
rect 132034 77568 132040 77580
rect 131724 77540 132040 77568
rect 131724 77528 131730 77540
rect 132034 77528 132040 77540
rect 132092 77528 132098 77580
rect 136634 77528 136640 77580
rect 136692 77568 136698 77580
rect 139026 77568 139032 77580
rect 136692 77540 139032 77568
rect 136692 77528 136698 77540
rect 139026 77528 139032 77540
rect 139084 77528 139090 77580
rect 130010 77460 130016 77512
rect 130068 77500 130074 77512
rect 135622 77500 135628 77512
rect 130068 77472 135628 77500
rect 130068 77460 130074 77472
rect 135622 77460 135628 77472
rect 135680 77460 135686 77512
rect 147766 77460 147772 77512
rect 147824 77500 147830 77512
rect 154684 77500 154712 77676
rect 158346 77664 158352 77716
rect 158404 77704 158410 77716
rect 172422 77704 172428 77716
rect 158404 77676 172428 77704
rect 158404 77664 158410 77676
rect 172422 77664 172428 77676
rect 172480 77664 172486 77716
rect 159910 77596 159916 77648
rect 159968 77636 159974 77648
rect 171410 77636 171416 77648
rect 159968 77608 171416 77636
rect 159968 77596 159974 77608
rect 171410 77596 171416 77608
rect 171468 77596 171474 77648
rect 160370 77528 160376 77580
rect 160428 77568 160434 77580
rect 160646 77568 160652 77580
rect 160428 77540 160652 77568
rect 160428 77528 160434 77540
rect 160646 77528 160652 77540
rect 160704 77528 160710 77580
rect 171594 77528 171600 77580
rect 171652 77568 171658 77580
rect 580626 77568 580632 77580
rect 171652 77540 580632 77568
rect 171652 77528 171658 77540
rect 580626 77528 580632 77540
rect 580684 77528 580690 77580
rect 167454 77500 167460 77512
rect 147824 77472 154574 77500
rect 154684 77472 167460 77500
rect 147824 77460 147830 77472
rect 126330 77392 126336 77444
rect 126388 77432 126394 77444
rect 130378 77432 130384 77444
rect 126388 77404 130384 77432
rect 126388 77392 126394 77404
rect 130378 77392 130384 77404
rect 130436 77392 130442 77444
rect 133506 77392 133512 77444
rect 133564 77432 133570 77444
rect 136910 77432 136916 77444
rect 133564 77404 136916 77432
rect 133564 77392 133570 77404
rect 136910 77392 136916 77404
rect 136968 77392 136974 77444
rect 149698 77392 149704 77444
rect 149756 77432 149762 77444
rect 152642 77432 152648 77444
rect 149756 77404 152648 77432
rect 149756 77392 149762 77404
rect 152642 77392 152648 77404
rect 152700 77392 152706 77444
rect 154546 77432 154574 77472
rect 167454 77460 167460 77472
rect 167512 77460 167518 77512
rect 168282 77460 168288 77512
rect 168340 77500 168346 77512
rect 171778 77500 171784 77512
rect 168340 77472 171784 77500
rect 168340 77460 168346 77472
rect 171778 77460 171784 77472
rect 171836 77460 171842 77512
rect 158254 77432 158260 77444
rect 154546 77404 158260 77432
rect 158254 77392 158260 77404
rect 158312 77392 158318 77444
rect 171318 77392 171324 77444
rect 171376 77432 171382 77444
rect 171686 77432 171692 77444
rect 171376 77404 171692 77432
rect 171376 77392 171382 77404
rect 171686 77392 171692 77404
rect 171744 77392 171750 77444
rect 144914 77324 144920 77376
rect 144972 77364 144978 77376
rect 162210 77364 162216 77376
rect 144972 77336 162216 77364
rect 144972 77324 144978 77336
rect 162210 77324 162216 77336
rect 162268 77324 162274 77376
rect 163406 77324 163412 77376
rect 163464 77364 163470 77376
rect 172054 77364 172060 77376
rect 163464 77336 172060 77364
rect 163464 77324 163470 77336
rect 172054 77324 172060 77336
rect 172112 77324 172118 77376
rect 142430 77256 142436 77308
rect 142488 77296 142494 77308
rect 142798 77296 142804 77308
rect 142488 77268 142804 77296
rect 142488 77256 142494 77268
rect 142798 77256 142804 77268
rect 142856 77256 142862 77308
rect 148870 77256 148876 77308
rect 148928 77296 148934 77308
rect 148928 77268 150434 77296
rect 148928 77256 148934 77268
rect 148962 77188 148968 77240
rect 149020 77228 149026 77240
rect 149514 77228 149520 77240
rect 149020 77200 149520 77228
rect 149020 77188 149026 77200
rect 149514 77188 149520 77200
rect 149572 77188 149578 77240
rect 150406 77228 150434 77268
rect 151262 77256 151268 77308
rect 151320 77296 151326 77308
rect 151320 77268 154252 77296
rect 151320 77256 151326 77268
rect 154224 77240 154252 77268
rect 156138 77256 156144 77308
rect 156196 77296 156202 77308
rect 157058 77296 157064 77308
rect 156196 77268 157064 77296
rect 156196 77256 156202 77268
rect 157058 77256 157064 77268
rect 157116 77256 157122 77308
rect 153010 77228 153016 77240
rect 150406 77200 153016 77228
rect 153010 77188 153016 77200
rect 153068 77188 153074 77240
rect 154206 77188 154212 77240
rect 154264 77188 154270 77240
rect 178770 77188 178776 77240
rect 178828 77228 178834 77240
rect 527174 77228 527180 77240
rect 178828 77200 527180 77228
rect 178828 77188 178834 77200
rect 527174 77188 527180 77200
rect 527232 77188 527238 77240
rect 120902 77120 120908 77172
rect 120960 77160 120966 77172
rect 171870 77160 171876 77172
rect 120960 77132 171876 77160
rect 120960 77120 120966 77132
rect 171870 77120 171876 77132
rect 171928 77120 171934 77172
rect 120994 77052 121000 77104
rect 121052 77092 121058 77104
rect 172606 77092 172612 77104
rect 121052 77064 172612 77092
rect 121052 77052 121058 77064
rect 172606 77052 172612 77064
rect 172664 77052 172670 77104
rect 153838 76984 153844 77036
rect 153896 77024 153902 77036
rect 211798 77024 211804 77036
rect 153896 76996 211804 77024
rect 153896 76984 153902 76996
rect 211798 76984 211804 76996
rect 211856 76984 211862 77036
rect 152366 76916 152372 76968
rect 152424 76956 152430 76968
rect 226334 76956 226340 76968
rect 152424 76928 226340 76956
rect 152424 76916 152430 76928
rect 226334 76916 226340 76928
rect 226392 76916 226398 76968
rect 124858 76848 124864 76900
rect 124916 76888 124922 76900
rect 134794 76888 134800 76900
rect 124916 76860 134800 76888
rect 124916 76848 124922 76860
rect 134794 76848 134800 76860
rect 134852 76848 134858 76900
rect 146938 76848 146944 76900
rect 146996 76888 147002 76900
rect 240134 76888 240140 76900
rect 146996 76860 240140 76888
rect 146996 76848 147002 76860
rect 240134 76848 240140 76860
rect 240192 76848 240198 76900
rect 102134 76780 102140 76832
rect 102192 76820 102198 76832
rect 132494 76820 132500 76832
rect 102192 76792 132500 76820
rect 102192 76780 102198 76792
rect 132494 76780 132500 76792
rect 132552 76780 132558 76832
rect 135622 76780 135628 76832
rect 135680 76820 135686 76832
rect 135806 76820 135812 76832
rect 135680 76792 135812 76820
rect 135680 76780 135686 76792
rect 135806 76780 135812 76792
rect 135864 76780 135870 76832
rect 145650 76780 145656 76832
rect 145708 76820 145714 76832
rect 260834 76820 260840 76832
rect 145708 76792 260840 76820
rect 145708 76780 145714 76792
rect 260834 76780 260840 76792
rect 260892 76780 260898 76832
rect 86954 76712 86960 76764
rect 87012 76752 87018 76764
rect 132310 76752 132316 76764
rect 87012 76724 132316 76752
rect 87012 76712 87018 76724
rect 132310 76712 132316 76724
rect 132368 76712 132374 76764
rect 148318 76712 148324 76764
rect 148376 76752 148382 76764
rect 148376 76724 152826 76752
rect 148376 76712 148382 76724
rect 69014 76644 69020 76696
rect 69072 76684 69078 76696
rect 128538 76684 128544 76696
rect 69072 76656 128544 76684
rect 69072 76644 69078 76656
rect 128538 76644 128544 76656
rect 128596 76644 128602 76696
rect 132586 76644 132592 76696
rect 132644 76684 132650 76696
rect 133138 76684 133144 76696
rect 132644 76656 133144 76684
rect 132644 76644 132650 76656
rect 133138 76644 133144 76656
rect 133196 76644 133202 76696
rect 145466 76644 145472 76696
rect 145524 76684 145530 76696
rect 145650 76684 145656 76696
rect 145524 76656 145656 76684
rect 145524 76644 145530 76656
rect 145650 76644 145656 76656
rect 145708 76644 145714 76696
rect 150526 76644 150532 76696
rect 150584 76684 150590 76696
rect 152798 76684 152826 76724
rect 153010 76712 153016 76764
rect 153068 76752 153074 76764
rect 288434 76752 288440 76764
rect 153068 76724 288440 76752
rect 153068 76712 153074 76724
rect 288434 76712 288440 76724
rect 288492 76712 288498 76764
rect 296714 76684 296720 76696
rect 150584 76656 152504 76684
rect 152798 76656 296720 76684
rect 150584 76644 150590 76656
rect 44174 76576 44180 76628
rect 44232 76616 44238 76628
rect 128354 76616 128360 76628
rect 44232 76588 128360 76616
rect 44232 76576 44238 76588
rect 128354 76576 128360 76588
rect 128412 76576 128418 76628
rect 143166 76576 143172 76628
rect 143224 76616 143230 76628
rect 152366 76616 152372 76628
rect 143224 76588 152372 76616
rect 143224 76576 143230 76588
rect 152366 76576 152372 76588
rect 152424 76576 152430 76628
rect 152476 76616 152504 76656
rect 296714 76644 296720 76656
rect 296772 76644 296778 76696
rect 324406 76616 324412 76628
rect 152476 76588 324412 76616
rect 324406 76576 324412 76588
rect 324464 76576 324470 76628
rect 30374 76508 30380 76560
rect 30432 76548 30438 76560
rect 127894 76548 127900 76560
rect 30432 76520 127900 76548
rect 30432 76508 30438 76520
rect 127894 76508 127900 76520
rect 127952 76508 127958 76560
rect 137370 76508 137376 76560
rect 137428 76548 137434 76560
rect 144546 76548 144552 76560
rect 137428 76520 144552 76548
rect 137428 76508 137434 76520
rect 144546 76508 144552 76520
rect 144604 76508 144610 76560
rect 152090 76508 152096 76560
rect 152148 76548 152154 76560
rect 152274 76548 152280 76560
rect 152148 76520 152280 76548
rect 152148 76508 152154 76520
rect 152274 76508 152280 76520
rect 152332 76508 152338 76560
rect 158714 76508 158720 76560
rect 158772 76548 158778 76560
rect 159266 76548 159272 76560
rect 158772 76520 159272 76548
rect 158772 76508 158778 76520
rect 159266 76508 159272 76520
rect 159324 76508 159330 76560
rect 159450 76508 159456 76560
rect 159508 76548 159514 76560
rect 160002 76548 160008 76560
rect 159508 76520 160008 76548
rect 159508 76508 159514 76520
rect 160002 76508 160008 76520
rect 160060 76508 160066 76560
rect 160186 76508 160192 76560
rect 160244 76548 160250 76560
rect 454034 76548 454040 76560
rect 160244 76520 454040 76548
rect 160244 76508 160250 76520
rect 454034 76508 454040 76520
rect 454092 76508 454098 76560
rect 122834 76440 122840 76492
rect 122892 76480 122898 76492
rect 135070 76480 135076 76492
rect 122892 76452 135076 76480
rect 122892 76440 122898 76452
rect 135070 76440 135076 76452
rect 135128 76440 135134 76492
rect 150250 76440 150256 76492
rect 150308 76480 150314 76492
rect 197354 76480 197360 76492
rect 150308 76452 197360 76480
rect 150308 76440 150314 76452
rect 197354 76440 197360 76452
rect 197412 76440 197418 76492
rect 119982 76372 119988 76424
rect 120040 76412 120046 76424
rect 172882 76412 172888 76424
rect 120040 76384 172888 76412
rect 120040 76372 120046 76384
rect 172882 76372 172888 76384
rect 172940 76372 172946 76424
rect 127618 76304 127624 76356
rect 127676 76344 127682 76356
rect 129182 76344 129188 76356
rect 127676 76316 129188 76344
rect 127676 76304 127682 76316
rect 129182 76304 129188 76316
rect 129240 76304 129246 76356
rect 156046 76304 156052 76356
rect 156104 76344 156110 76356
rect 156414 76344 156420 76356
rect 156104 76316 156420 76344
rect 156104 76304 156110 76316
rect 156414 76304 156420 76316
rect 156472 76304 156478 76356
rect 158714 76304 158720 76356
rect 158772 76344 158778 76356
rect 159726 76344 159732 76356
rect 158772 76316 159732 76344
rect 158772 76304 158778 76316
rect 159726 76304 159732 76316
rect 159784 76304 159790 76356
rect 127250 76236 127256 76288
rect 127308 76276 127314 76288
rect 128262 76276 128268 76288
rect 127308 76248 128268 76276
rect 127308 76236 127314 76248
rect 128262 76236 128268 76248
rect 128320 76236 128326 76288
rect 151814 76236 151820 76288
rect 151872 76276 151878 76288
rect 152274 76276 152280 76288
rect 151872 76248 152280 76276
rect 151872 76236 151878 76248
rect 152274 76236 152280 76248
rect 152332 76236 152338 76288
rect 155770 76236 155776 76288
rect 155828 76276 155834 76288
rect 159634 76276 159640 76288
rect 155828 76248 159640 76276
rect 155828 76236 155834 76248
rect 159634 76236 159640 76248
rect 159692 76236 159698 76288
rect 143626 76168 143632 76220
rect 143684 76208 143690 76220
rect 144086 76208 144092 76220
rect 143684 76180 144092 76208
rect 143684 76168 143690 76180
rect 144086 76168 144092 76180
rect 144144 76168 144150 76220
rect 154574 76168 154580 76220
rect 154632 76208 154638 76220
rect 155126 76208 155132 76220
rect 154632 76180 155132 76208
rect 154632 76168 154638 76180
rect 155126 76168 155132 76180
rect 155184 76168 155190 76220
rect 154666 76100 154672 76152
rect 154724 76140 154730 76152
rect 155218 76140 155224 76152
rect 154724 76112 155224 76140
rect 154724 76100 154730 76112
rect 155218 76100 155224 76112
rect 155276 76100 155282 76152
rect 143810 76032 143816 76084
rect 143868 76032 143874 76084
rect 143902 76032 143908 76084
rect 143960 76072 143966 76084
rect 144086 76072 144092 76084
rect 143960 76044 144092 76072
rect 143960 76032 143966 76044
rect 144086 76032 144092 76044
rect 144144 76032 144150 76084
rect 153470 76032 153476 76084
rect 153528 76072 153534 76084
rect 155862 76072 155868 76084
rect 153528 76044 155868 76072
rect 153528 76032 153534 76044
rect 155862 76032 155868 76044
rect 155920 76032 155926 76084
rect 156230 76032 156236 76084
rect 156288 76072 156294 76084
rect 156506 76072 156512 76084
rect 156288 76044 156512 76072
rect 156288 76032 156294 76044
rect 156506 76032 156512 76044
rect 156564 76032 156570 76084
rect 125502 75896 125508 75948
rect 125560 75936 125566 75948
rect 126238 75936 126244 75948
rect 125560 75908 126244 75936
rect 125560 75896 125566 75908
rect 126238 75896 126244 75908
rect 126296 75896 126302 75948
rect 127434 75896 127440 75948
rect 127492 75936 127498 75948
rect 127710 75936 127716 75948
rect 127492 75908 127716 75936
rect 127492 75896 127498 75908
rect 127710 75896 127716 75908
rect 127768 75896 127774 75948
rect 141050 75896 141056 75948
rect 141108 75936 141114 75948
rect 141694 75936 141700 75948
rect 141108 75908 141700 75936
rect 141108 75896 141114 75908
rect 141694 75896 141700 75908
rect 141752 75896 141758 75948
rect 142154 75896 142160 75948
rect 142212 75936 142218 75948
rect 143074 75936 143080 75948
rect 142212 75908 143080 75936
rect 142212 75896 142218 75908
rect 143074 75896 143080 75908
rect 143132 75896 143138 75948
rect 143828 75936 143856 76032
rect 143902 75936 143908 75948
rect 143828 75908 143908 75936
rect 143902 75896 143908 75908
rect 143960 75896 143966 75948
rect 153378 75896 153384 75948
rect 153436 75936 153442 75948
rect 154114 75936 154120 75948
rect 153436 75908 154120 75936
rect 153436 75896 153442 75908
rect 154114 75896 154120 75908
rect 154172 75896 154178 75948
rect 154574 75896 154580 75948
rect 154632 75936 154638 75948
rect 155494 75936 155500 75948
rect 154632 75908 155500 75936
rect 154632 75896 154638 75908
rect 155494 75896 155500 75908
rect 155552 75896 155558 75948
rect 157242 75896 157248 75948
rect 157300 75936 157306 75948
rect 158254 75936 158260 75948
rect 157300 75908 158260 75936
rect 157300 75896 157306 75908
rect 158254 75896 158260 75908
rect 158312 75896 158318 75948
rect 122098 75828 122104 75880
rect 122156 75868 122162 75880
rect 127342 75868 127348 75880
rect 122156 75840 127348 75868
rect 122156 75828 122162 75840
rect 127342 75828 127348 75840
rect 127400 75828 127406 75880
rect 153286 75828 153292 75880
rect 153344 75868 153350 75880
rect 153562 75868 153568 75880
rect 153344 75840 153568 75868
rect 153344 75828 153350 75840
rect 153562 75828 153568 75840
rect 153620 75828 153626 75880
rect 155954 75828 155960 75880
rect 156012 75868 156018 75880
rect 156598 75868 156604 75880
rect 156012 75840 156604 75868
rect 156012 75828 156018 75840
rect 156598 75828 156604 75840
rect 156656 75828 156662 75880
rect 120718 75760 120724 75812
rect 120776 75800 120782 75812
rect 128446 75800 128452 75812
rect 120776 75772 128452 75800
rect 120776 75760 120782 75772
rect 128446 75760 128452 75772
rect 128504 75760 128510 75812
rect 154758 75760 154764 75812
rect 154816 75800 154822 75812
rect 155034 75800 155040 75812
rect 154816 75772 155040 75800
rect 154816 75760 154822 75772
rect 155034 75760 155040 75772
rect 155092 75760 155098 75812
rect 156782 75760 156788 75812
rect 156840 75800 156846 75812
rect 156840 75772 173894 75800
rect 156840 75760 156846 75772
rect 127342 75692 127348 75744
rect 127400 75732 127406 75744
rect 128170 75732 128176 75744
rect 127400 75704 128176 75732
rect 127400 75692 127406 75704
rect 128170 75692 128176 75704
rect 128228 75692 128234 75744
rect 129826 75692 129832 75744
rect 129884 75732 129890 75744
rect 130010 75732 130016 75744
rect 129884 75704 130016 75732
rect 129884 75692 129890 75704
rect 130010 75692 130016 75704
rect 130068 75692 130074 75744
rect 142246 75692 142252 75744
rect 142304 75732 142310 75744
rect 142982 75732 142988 75744
rect 142304 75704 142988 75732
rect 142304 75692 142310 75704
rect 142982 75692 142988 75704
rect 143040 75692 143046 75744
rect 151814 75692 151820 75744
rect 151872 75732 151878 75744
rect 152182 75732 152188 75744
rect 151872 75704 152188 75732
rect 151872 75692 151878 75704
rect 152182 75692 152188 75704
rect 152240 75692 152246 75744
rect 122282 75624 122288 75676
rect 122340 75664 122346 75676
rect 128078 75664 128084 75676
rect 122340 75636 128084 75664
rect 122340 75624 122346 75636
rect 128078 75624 128084 75636
rect 128136 75624 128142 75676
rect 158990 75624 158996 75676
rect 159048 75664 159054 75676
rect 159048 75636 166994 75664
rect 159048 75624 159054 75636
rect 130010 75556 130016 75608
rect 130068 75596 130074 75608
rect 130654 75596 130660 75608
rect 130068 75568 130660 75596
rect 130068 75556 130074 75568
rect 130654 75556 130660 75568
rect 130712 75556 130718 75608
rect 159910 75556 159916 75608
rect 159968 75596 159974 75608
rect 166718 75596 166724 75608
rect 159968 75568 166724 75596
rect 159968 75556 159974 75568
rect 166718 75556 166724 75568
rect 166776 75556 166782 75608
rect 122190 75488 122196 75540
rect 122248 75528 122254 75540
rect 130470 75528 130476 75540
rect 122248 75500 130476 75528
rect 122248 75488 122254 75500
rect 130470 75488 130476 75500
rect 130528 75488 130534 75540
rect 154758 75488 154764 75540
rect 154816 75528 154822 75540
rect 155402 75528 155408 75540
rect 154816 75500 155408 75528
rect 154816 75488 154822 75500
rect 155402 75488 155408 75500
rect 155460 75488 155466 75540
rect 162210 75488 162216 75540
rect 162268 75528 162274 75540
rect 166966 75528 166994 75636
rect 173866 75596 173894 75772
rect 396074 75596 396080 75608
rect 173866 75568 396080 75596
rect 396074 75556 396080 75568
rect 396132 75556 396138 75608
rect 431954 75528 431960 75540
rect 162268 75500 166764 75528
rect 166966 75500 431960 75528
rect 162268 75488 162274 75500
rect 121454 75420 121460 75472
rect 121512 75460 121518 75472
rect 134978 75460 134984 75472
rect 121512 75432 134984 75460
rect 121512 75420 121518 75432
rect 134978 75420 134984 75432
rect 135036 75420 135042 75472
rect 136818 75420 136824 75472
rect 136876 75460 136882 75472
rect 137646 75460 137652 75472
rect 136876 75432 137652 75460
rect 136876 75420 136882 75432
rect 137646 75420 137652 75432
rect 137704 75420 137710 75472
rect 163958 75420 163964 75472
rect 164016 75460 164022 75472
rect 164016 75432 166672 75460
rect 164016 75420 164022 75432
rect 51074 75352 51080 75404
rect 51132 75392 51138 75404
rect 129090 75392 129096 75404
rect 51132 75364 129096 75392
rect 51132 75352 51138 75364
rect 129090 75352 129096 75364
rect 129148 75352 129154 75404
rect 136910 75352 136916 75404
rect 136968 75392 136974 75404
rect 137278 75392 137284 75404
rect 136968 75364 137284 75392
rect 136968 75352 136974 75364
rect 137278 75352 137284 75364
rect 137336 75352 137342 75404
rect 149330 75352 149336 75404
rect 149388 75392 149394 75404
rect 149514 75392 149520 75404
rect 149388 75364 149520 75392
rect 149388 75352 149394 75364
rect 149514 75352 149520 75364
rect 149572 75352 149578 75404
rect 155954 75352 155960 75404
rect 156012 75392 156018 75404
rect 156690 75392 156696 75404
rect 156012 75364 156696 75392
rect 156012 75352 156018 75364
rect 156690 75352 156696 75364
rect 156748 75352 156754 75404
rect 164418 75352 164424 75404
rect 164476 75392 164482 75404
rect 164694 75392 164700 75404
rect 164476 75364 164700 75392
rect 164476 75352 164482 75364
rect 164694 75352 164700 75364
rect 164752 75352 164758 75404
rect 165798 75352 165804 75404
rect 165856 75392 165862 75404
rect 166534 75392 166540 75404
rect 165856 75364 166540 75392
rect 165856 75352 165862 75364
rect 166534 75352 166540 75364
rect 166592 75352 166598 75404
rect 107654 75284 107660 75336
rect 107712 75324 107718 75336
rect 131574 75324 131580 75336
rect 107712 75296 131580 75324
rect 107712 75284 107718 75296
rect 131574 75284 131580 75296
rect 131632 75284 131638 75336
rect 132678 75284 132684 75336
rect 132736 75324 132742 75336
rect 133598 75324 133604 75336
rect 132736 75296 133604 75324
rect 132736 75284 132742 75296
rect 133598 75284 133604 75296
rect 133656 75284 133662 75336
rect 135438 75284 135444 75336
rect 135496 75324 135502 75336
rect 136174 75324 136180 75336
rect 135496 75296 136180 75324
rect 135496 75284 135502 75296
rect 136174 75284 136180 75296
rect 136232 75284 136238 75336
rect 144914 75284 144920 75336
rect 144972 75324 144978 75336
rect 145834 75324 145840 75336
rect 144972 75296 145840 75324
rect 144972 75284 144978 75296
rect 145834 75284 145840 75296
rect 145892 75284 145898 75336
rect 146202 75284 146208 75336
rect 146260 75324 146266 75336
rect 146846 75324 146852 75336
rect 146260 75296 146852 75324
rect 146260 75284 146266 75296
rect 146846 75284 146852 75296
rect 146904 75284 146910 75336
rect 147674 75284 147680 75336
rect 147732 75324 147738 75336
rect 148594 75324 148600 75336
rect 147732 75296 148600 75324
rect 147732 75284 147738 75296
rect 148594 75284 148600 75296
rect 148652 75284 148658 75336
rect 151906 75284 151912 75336
rect 151964 75324 151970 75336
rect 152366 75324 152372 75336
rect 151964 75296 152372 75324
rect 151964 75284 151970 75296
rect 152366 75284 152372 75296
rect 152424 75284 152430 75336
rect 164602 75284 164608 75336
rect 164660 75324 164666 75336
rect 166644 75324 166672 75432
rect 166736 75392 166764 75500
rect 431954 75488 431960 75500
rect 432012 75488 432018 75540
rect 166810 75420 166816 75472
rect 166868 75460 166874 75472
rect 438854 75460 438860 75472
rect 166868 75432 438860 75460
rect 166868 75420 166874 75432
rect 438854 75420 438860 75432
rect 438912 75420 438918 75472
rect 467834 75392 467840 75404
rect 166736 75364 467840 75392
rect 467834 75352 467840 75364
rect 467892 75352 467898 75404
rect 490006 75324 490012 75336
rect 164660 75296 166488 75324
rect 166644 75296 490012 75324
rect 164660 75284 164666 75296
rect 42794 75216 42800 75268
rect 42852 75256 42858 75268
rect 128354 75256 128360 75268
rect 42852 75228 128360 75256
rect 42852 75216 42858 75228
rect 128354 75216 128360 75228
rect 128412 75216 128418 75268
rect 128722 75216 128728 75268
rect 128780 75256 128786 75268
rect 129642 75256 129648 75268
rect 128780 75228 129648 75256
rect 128780 75216 128786 75228
rect 129642 75216 129648 75228
rect 129700 75216 129706 75268
rect 130286 75216 130292 75268
rect 130344 75256 130350 75268
rect 131022 75256 131028 75268
rect 130344 75228 131028 75256
rect 130344 75216 130350 75228
rect 131022 75216 131028 75228
rect 131080 75216 131086 75268
rect 132862 75216 132868 75268
rect 132920 75256 132926 75268
rect 133690 75256 133696 75268
rect 132920 75228 133696 75256
rect 132920 75216 132926 75228
rect 133690 75216 133696 75228
rect 133748 75216 133754 75268
rect 134242 75216 134248 75268
rect 134300 75256 134306 75268
rect 134702 75256 134708 75268
rect 134300 75228 134708 75256
rect 134300 75216 134306 75228
rect 134702 75216 134708 75228
rect 134760 75216 134766 75268
rect 135898 75216 135904 75268
rect 135956 75256 135962 75268
rect 136358 75256 136364 75268
rect 135956 75228 136364 75256
rect 135956 75216 135962 75228
rect 136358 75216 136364 75228
rect 136416 75216 136422 75268
rect 136818 75216 136824 75268
rect 136876 75256 136882 75268
rect 137462 75256 137468 75268
rect 136876 75228 137468 75256
rect 136876 75216 136882 75228
rect 137462 75216 137468 75228
rect 137520 75216 137526 75268
rect 138106 75216 138112 75268
rect 138164 75256 138170 75268
rect 138658 75256 138664 75268
rect 138164 75228 138664 75256
rect 138164 75216 138170 75228
rect 138658 75216 138664 75228
rect 138716 75216 138722 75268
rect 139670 75216 139676 75268
rect 139728 75256 139734 75268
rect 140130 75256 140136 75268
rect 139728 75228 140136 75256
rect 139728 75216 139734 75228
rect 140130 75216 140136 75228
rect 140188 75216 140194 75268
rect 143994 75216 144000 75268
rect 144052 75256 144058 75268
rect 144454 75256 144460 75268
rect 144052 75228 144460 75256
rect 144052 75216 144058 75228
rect 144454 75216 144460 75228
rect 144512 75216 144518 75268
rect 145374 75216 145380 75268
rect 145432 75256 145438 75268
rect 145742 75256 145748 75268
rect 145432 75228 145748 75256
rect 145432 75216 145438 75228
rect 145742 75216 145748 75228
rect 145800 75216 145806 75268
rect 146478 75216 146484 75268
rect 146536 75256 146542 75268
rect 146754 75256 146760 75268
rect 146536 75228 146760 75256
rect 146536 75216 146542 75228
rect 146754 75216 146760 75228
rect 146812 75216 146818 75268
rect 146938 75216 146944 75268
rect 146996 75256 147002 75268
rect 147122 75256 147128 75268
rect 146996 75228 147128 75256
rect 146996 75216 147002 75228
rect 147122 75216 147128 75228
rect 147180 75216 147186 75268
rect 148042 75216 148048 75268
rect 148100 75256 148106 75268
rect 148410 75256 148416 75268
rect 148100 75228 148416 75256
rect 148100 75216 148106 75228
rect 148410 75216 148416 75228
rect 148468 75216 148474 75268
rect 149330 75216 149336 75268
rect 149388 75256 149394 75268
rect 149882 75256 149888 75268
rect 149388 75228 149888 75256
rect 149388 75216 149394 75228
rect 149882 75216 149888 75228
rect 149940 75216 149946 75268
rect 150710 75216 150716 75268
rect 150768 75256 150774 75268
rect 151078 75256 151084 75268
rect 150768 75228 151084 75256
rect 150768 75216 150774 75228
rect 151078 75216 151084 75228
rect 151136 75216 151142 75268
rect 152182 75216 152188 75268
rect 152240 75256 152246 75268
rect 152550 75256 152556 75268
rect 152240 75228 152556 75256
rect 152240 75216 152246 75228
rect 152550 75216 152556 75228
rect 152608 75216 152614 75268
rect 153194 75216 153200 75268
rect 153252 75256 153258 75268
rect 153930 75256 153936 75268
rect 153252 75228 153936 75256
rect 153252 75216 153258 75228
rect 153930 75216 153936 75228
rect 153988 75216 153994 75268
rect 157518 75216 157524 75268
rect 157576 75256 157582 75268
rect 158070 75256 158076 75268
rect 157576 75228 158076 75256
rect 157576 75216 157582 75228
rect 158070 75216 158076 75228
rect 158128 75216 158134 75268
rect 160370 75216 160376 75268
rect 160428 75256 160434 75268
rect 160738 75256 160744 75268
rect 160428 75228 160744 75256
rect 160428 75216 160434 75228
rect 160738 75216 160744 75228
rect 160796 75216 160802 75268
rect 161566 75216 161572 75268
rect 161624 75256 161630 75268
rect 162026 75256 162032 75268
rect 161624 75228 162032 75256
rect 161624 75216 161630 75228
rect 162026 75216 162032 75228
rect 162084 75216 162090 75268
rect 163038 75216 163044 75268
rect 163096 75256 163102 75268
rect 163406 75256 163412 75268
rect 163096 75228 163412 75256
rect 163096 75216 163102 75228
rect 163406 75216 163412 75228
rect 163464 75216 163470 75268
rect 164694 75216 164700 75268
rect 164752 75256 164758 75268
rect 164970 75256 164976 75268
rect 164752 75228 164976 75256
rect 164752 75216 164758 75228
rect 164970 75216 164976 75228
rect 165028 75216 165034 75268
rect 165798 75216 165804 75268
rect 165856 75256 165862 75268
rect 166350 75256 166356 75268
rect 165856 75228 166356 75256
rect 165856 75216 165862 75228
rect 166350 75216 166356 75228
rect 166408 75216 166414 75268
rect 166460 75256 166488 75296
rect 490006 75284 490012 75296
rect 490064 75284 490070 75336
rect 499574 75256 499580 75268
rect 166460 75228 499580 75256
rect 499574 75216 499580 75228
rect 499632 75216 499638 75268
rect 6914 75148 6920 75200
rect 6972 75188 6978 75200
rect 123018 75188 123024 75200
rect 6972 75160 123024 75188
rect 6972 75148 6978 75160
rect 123018 75148 123024 75160
rect 123076 75148 123082 75200
rect 128538 75148 128544 75200
rect 128596 75188 128602 75200
rect 128906 75188 128912 75200
rect 128596 75160 128912 75188
rect 128596 75148 128602 75160
rect 128906 75148 128912 75160
rect 128964 75148 128970 75200
rect 132954 75148 132960 75200
rect 133012 75188 133018 75200
rect 133782 75188 133788 75200
rect 133012 75160 133788 75188
rect 133012 75148 133018 75160
rect 133782 75148 133788 75160
rect 133840 75148 133846 75200
rect 135530 75148 135536 75200
rect 135588 75188 135594 75200
rect 136266 75188 136272 75200
rect 135588 75160 136272 75188
rect 135588 75148 135594 75160
rect 136266 75148 136272 75160
rect 136324 75148 136330 75200
rect 137002 75148 137008 75200
rect 137060 75188 137066 75200
rect 137186 75188 137192 75200
rect 137060 75160 137192 75188
rect 137060 75148 137066 75160
rect 137186 75148 137192 75160
rect 137244 75148 137250 75200
rect 139946 75148 139952 75200
rect 140004 75188 140010 75200
rect 140222 75188 140228 75200
rect 140004 75160 140228 75188
rect 140004 75148 140010 75160
rect 140222 75148 140228 75160
rect 140280 75148 140286 75200
rect 145098 75148 145104 75200
rect 145156 75188 145162 75200
rect 145466 75188 145472 75200
rect 145156 75160 145472 75188
rect 145156 75148 145162 75160
rect 145466 75148 145472 75160
rect 145524 75148 145530 75200
rect 146570 75148 146576 75200
rect 146628 75188 146634 75200
rect 146846 75188 146852 75200
rect 146628 75160 146852 75188
rect 146628 75148 146634 75160
rect 146846 75148 146852 75160
rect 146904 75148 146910 75200
rect 147766 75148 147772 75200
rect 147824 75188 147830 75200
rect 148502 75188 148508 75200
rect 147824 75160 148508 75188
rect 147824 75148 147830 75160
rect 148502 75148 148508 75160
rect 148560 75148 148566 75200
rect 151906 75148 151912 75200
rect 151964 75188 151970 75200
rect 152918 75188 152924 75200
rect 151964 75160 152924 75188
rect 151964 75148 151970 75160
rect 152918 75148 152924 75160
rect 152976 75148 152982 75200
rect 157794 75148 157800 75200
rect 157852 75188 157858 75200
rect 158162 75188 158168 75200
rect 157852 75160 158168 75188
rect 157852 75148 157858 75160
rect 158162 75148 158168 75160
rect 158220 75148 158226 75200
rect 160186 75148 160192 75200
rect 160244 75188 160250 75200
rect 160830 75188 160836 75200
rect 160244 75160 160836 75188
rect 160244 75148 160250 75160
rect 160830 75148 160836 75160
rect 160888 75148 160894 75200
rect 162854 75148 162860 75200
rect 162912 75188 162918 75200
rect 163498 75188 163504 75200
rect 162912 75160 163504 75188
rect 162912 75148 162918 75160
rect 163498 75148 163504 75160
rect 163556 75148 163562 75200
rect 164602 75148 164608 75200
rect 164660 75188 164666 75200
rect 165154 75188 165160 75200
rect 164660 75160 165160 75188
rect 164660 75148 164666 75160
rect 165154 75148 165160 75160
rect 165212 75148 165218 75200
rect 167454 75148 167460 75200
rect 167512 75188 167518 75200
rect 167822 75188 167828 75200
rect 167512 75160 167828 75188
rect 167512 75148 167518 75160
rect 167822 75148 167828 75160
rect 167880 75148 167886 75200
rect 168374 75148 168380 75200
rect 168432 75188 168438 75200
rect 168742 75188 168748 75200
rect 168432 75160 168748 75188
rect 168432 75148 168438 75160
rect 168742 75148 168748 75160
rect 168800 75148 168806 75200
rect 168834 75148 168840 75200
rect 168892 75188 168898 75200
rect 169386 75188 169392 75200
rect 168892 75160 169392 75188
rect 168892 75148 168898 75160
rect 169386 75148 169392 75160
rect 169444 75148 169450 75200
rect 169754 75148 169760 75200
rect 169812 75188 169818 75200
rect 170306 75188 170312 75200
rect 169812 75160 170312 75188
rect 169812 75148 169818 75160
rect 170306 75148 170312 75160
rect 170364 75148 170370 75200
rect 173986 75148 173992 75200
rect 174044 75188 174050 75200
rect 174354 75188 174360 75200
rect 174044 75160 174360 75188
rect 174044 75148 174050 75160
rect 174354 75148 174360 75160
rect 174412 75148 174418 75200
rect 564434 75188 564440 75200
rect 176626 75160 564440 75188
rect 128630 75080 128636 75132
rect 128688 75120 128694 75132
rect 129274 75120 129280 75132
rect 128688 75092 129280 75120
rect 128688 75080 128694 75092
rect 129274 75080 129280 75092
rect 129332 75080 129338 75132
rect 135714 75080 135720 75132
rect 135772 75120 135778 75132
rect 136450 75120 136456 75132
rect 135772 75092 136456 75120
rect 135772 75080 135778 75092
rect 136450 75080 136456 75092
rect 136508 75080 136514 75132
rect 138750 75080 138756 75132
rect 138808 75120 138814 75132
rect 140406 75120 140412 75132
rect 138808 75092 140412 75120
rect 138808 75080 138814 75092
rect 140406 75080 140412 75092
rect 140464 75080 140470 75132
rect 141234 75080 141240 75132
rect 141292 75120 141298 75132
rect 141510 75120 141516 75132
rect 141292 75092 141516 75120
rect 141292 75080 141298 75092
rect 141510 75080 141516 75092
rect 141568 75080 141574 75132
rect 142522 75080 142528 75132
rect 142580 75120 142586 75132
rect 142798 75120 142804 75132
rect 142580 75092 142804 75120
rect 142580 75080 142586 75092
rect 142798 75080 142804 75092
rect 142856 75080 142862 75132
rect 146478 75080 146484 75132
rect 146536 75120 146542 75132
rect 147490 75120 147496 75132
rect 146536 75092 147496 75120
rect 146536 75080 146542 75092
rect 147490 75080 147496 75092
rect 147548 75080 147554 75132
rect 150710 75080 150716 75132
rect 150768 75120 150774 75132
rect 151354 75120 151360 75132
rect 150768 75092 151360 75120
rect 150768 75080 150774 75092
rect 151354 75080 151360 75092
rect 151412 75080 151418 75132
rect 161566 75080 161572 75132
rect 161624 75120 161630 75132
rect 162118 75120 162124 75132
rect 161624 75092 162124 75120
rect 161624 75080 161630 75092
rect 162118 75080 162124 75092
rect 162176 75080 162182 75132
rect 163038 75080 163044 75132
rect 163096 75120 163102 75132
rect 163866 75120 163872 75132
rect 163096 75092 163872 75120
rect 163096 75080 163102 75092
rect 163866 75080 163872 75092
rect 163924 75080 163930 75132
rect 167086 75080 167092 75132
rect 167144 75120 167150 75132
rect 167914 75120 167920 75132
rect 167144 75092 167920 75120
rect 167144 75080 167150 75092
rect 167914 75080 167920 75092
rect 167972 75080 167978 75132
rect 170214 75080 170220 75132
rect 170272 75120 170278 75132
rect 170858 75120 170864 75132
rect 170272 75092 170864 75120
rect 170272 75080 170278 75092
rect 170858 75080 170864 75092
rect 170916 75080 170922 75132
rect 128354 75012 128360 75064
rect 128412 75052 128418 75064
rect 136542 75052 136548 75064
rect 128412 75024 136548 75052
rect 128412 75012 128418 75024
rect 136542 75012 136548 75024
rect 136600 75012 136606 75064
rect 137002 75012 137008 75064
rect 137060 75052 137066 75064
rect 137738 75052 137744 75064
rect 137060 75024 137744 75052
rect 137060 75012 137066 75024
rect 137738 75012 137744 75024
rect 137796 75012 137802 75064
rect 145098 75012 145104 75064
rect 145156 75052 145162 75064
rect 145926 75052 145932 75064
rect 145156 75024 145932 75052
rect 145156 75012 145162 75024
rect 145926 75012 145932 75024
rect 145984 75012 145990 75064
rect 146570 75012 146576 75064
rect 146628 75052 146634 75064
rect 147214 75052 147220 75064
rect 146628 75024 147220 75052
rect 146628 75012 146634 75024
rect 147214 75012 147220 75024
rect 147272 75012 147278 75064
rect 168374 75012 168380 75064
rect 168432 75052 168438 75064
rect 168558 75052 168564 75064
rect 168432 75024 168564 75052
rect 168432 75012 168438 75024
rect 168558 75012 168564 75024
rect 168616 75012 168622 75064
rect 169754 75012 169760 75064
rect 169812 75052 169818 75064
rect 170490 75052 170496 75064
rect 169812 75024 170496 75052
rect 169812 75012 169818 75024
rect 170490 75012 170496 75024
rect 170548 75012 170554 75064
rect 140958 74944 140964 74996
rect 141016 74984 141022 74996
rect 141786 74984 141792 74996
rect 141016 74956 141792 74984
rect 141016 74944 141022 74956
rect 141786 74944 141792 74956
rect 141844 74944 141850 74996
rect 169570 74944 169576 74996
rect 169628 74984 169634 74996
rect 176626 74984 176654 75160
rect 564434 75148 564440 75160
rect 564492 75148 564498 75200
rect 169628 74956 176654 74984
rect 169628 74944 169634 74956
rect 131666 74876 131672 74928
rect 131724 74916 131730 74928
rect 132126 74916 132132 74928
rect 131724 74888 132132 74916
rect 131724 74876 131730 74888
rect 132126 74876 132132 74888
rect 132184 74876 132190 74928
rect 146294 74876 146300 74928
rect 146352 74916 146358 74928
rect 147214 74916 147220 74928
rect 146352 74888 147220 74916
rect 146352 74876 146358 74888
rect 147214 74876 147220 74888
rect 147272 74876 147278 74928
rect 168558 74876 168564 74928
rect 168616 74916 168622 74928
rect 169110 74916 169116 74928
rect 168616 74888 169116 74916
rect 168616 74876 168622 74888
rect 169110 74876 169116 74888
rect 169168 74876 169174 74928
rect 124766 74808 124772 74860
rect 124824 74848 124830 74860
rect 125410 74848 125416 74860
rect 124824 74820 125416 74848
rect 124824 74808 124830 74820
rect 125410 74808 125416 74820
rect 125468 74808 125474 74860
rect 166994 74468 167000 74520
rect 167052 74508 167058 74520
rect 173342 74508 173348 74520
rect 167052 74480 173348 74508
rect 167052 74468 167058 74480
rect 173342 74468 173348 74480
rect 173400 74468 173406 74520
rect 141970 74196 141976 74248
rect 142028 74236 142034 74248
rect 209774 74236 209780 74248
rect 142028 74208 209780 74236
rect 142028 74196 142034 74208
rect 209774 74196 209780 74208
rect 209832 74196 209838 74248
rect 144822 74128 144828 74180
rect 144880 74168 144886 74180
rect 216674 74168 216680 74180
rect 144880 74140 216680 74168
rect 144880 74128 144886 74140
rect 216674 74128 216680 74140
rect 216732 74128 216738 74180
rect 118694 74060 118700 74112
rect 118752 74100 118758 74112
rect 134058 74100 134064 74112
rect 118752 74072 134064 74100
rect 118752 74060 118758 74072
rect 134058 74060 134064 74072
rect 134116 74060 134122 74112
rect 143442 74060 143448 74112
rect 143500 74100 143506 74112
rect 223574 74100 223580 74112
rect 143500 74072 223580 74100
rect 143500 74060 143506 74072
rect 223574 74060 223580 74072
rect 223632 74060 223638 74112
rect 93946 73992 93952 74044
rect 94004 74032 94010 74044
rect 133230 74032 133236 74044
rect 94004 74004 133236 74032
rect 94004 73992 94010 74004
rect 133230 73992 133236 74004
rect 133288 73992 133294 74044
rect 145650 73992 145656 74044
rect 145708 74032 145714 74044
rect 251174 74032 251180 74044
rect 145708 74004 251180 74032
rect 145708 73992 145714 74004
rect 251174 73992 251180 74004
rect 251232 73992 251238 74044
rect 64874 73924 64880 73976
rect 64932 73964 64938 73976
rect 129734 73964 129740 73976
rect 64932 73936 129740 73964
rect 64932 73924 64938 73936
rect 129734 73924 129740 73936
rect 129792 73924 129798 73976
rect 152642 73924 152648 73976
rect 152700 73964 152706 73976
rect 318794 73964 318800 73976
rect 152700 73936 318800 73964
rect 152700 73924 152706 73936
rect 318794 73924 318800 73936
rect 318852 73924 318858 73976
rect 27614 73856 27620 73908
rect 27672 73896 27678 73908
rect 126882 73896 126888 73908
rect 27672 73868 126888 73896
rect 27672 73856 27678 73868
rect 126882 73856 126888 73868
rect 126940 73856 126946 73908
rect 153102 73856 153108 73908
rect 153160 73896 153166 73908
rect 354674 73896 354680 73908
rect 153160 73868 354680 73896
rect 153160 73856 153166 73868
rect 354674 73856 354680 73868
rect 354732 73856 354738 73908
rect 26234 73788 26240 73840
rect 26292 73828 26298 73840
rect 122558 73828 122564 73840
rect 26292 73800 122564 73828
rect 26292 73788 26298 73800
rect 122558 73788 122564 73800
rect 122616 73788 122622 73840
rect 161014 73788 161020 73840
rect 161072 73828 161078 73840
rect 375374 73828 375380 73840
rect 161072 73800 375380 73828
rect 161072 73788 161078 73800
rect 375374 73788 375380 73800
rect 375432 73788 375438 73840
rect 137554 73176 137560 73228
rect 137612 73216 137618 73228
rect 142982 73216 142988 73228
rect 137612 73188 142988 73216
rect 137612 73176 137618 73188
rect 142982 73176 142988 73188
rect 143040 73176 143046 73228
rect 170950 73108 170956 73160
rect 171008 73148 171014 73160
rect 580166 73148 580172 73160
rect 171008 73120 580172 73148
rect 171008 73108 171014 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 126422 72768 126428 72820
rect 126480 72808 126486 72820
rect 126790 72808 126796 72820
rect 126480 72780 126796 72808
rect 126480 72768 126486 72780
rect 126790 72768 126796 72780
rect 126848 72768 126854 72820
rect 140866 72700 140872 72752
rect 140924 72740 140930 72752
rect 141418 72740 141424 72752
rect 140924 72712 141424 72740
rect 140924 72700 140930 72712
rect 141418 72700 141424 72712
rect 141476 72700 141482 72752
rect 148962 72632 148968 72684
rect 149020 72672 149026 72684
rect 291194 72672 291200 72684
rect 149020 72644 291200 72672
rect 149020 72632 149026 72644
rect 291194 72632 291200 72644
rect 291252 72632 291258 72684
rect 149054 72564 149060 72616
rect 149112 72604 149118 72616
rect 311894 72604 311900 72616
rect 149112 72576 311900 72604
rect 149112 72564 149118 72576
rect 311894 72564 311900 72576
rect 311952 72564 311958 72616
rect 152734 72496 152740 72548
rect 152792 72536 152798 72548
rect 340874 72536 340880 72548
rect 152792 72508 340880 72536
rect 152792 72496 152798 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 155862 72428 155868 72480
rect 155920 72468 155926 72480
rect 357434 72468 357440 72480
rect 155920 72440 357440 72468
rect 155920 72428 155926 72440
rect 357434 72428 357440 72440
rect 357492 72428 357498 72480
rect 165062 72360 165068 72412
rect 165120 72400 165126 72412
rect 171870 72400 171876 72412
rect 165120 72372 171876 72400
rect 165120 72360 165126 72372
rect 171870 72360 171876 72372
rect 171928 72360 171934 72412
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 179598 71720 179604 71732
rect 3476 71692 179604 71720
rect 3476 71680 3482 71692
rect 179598 71680 179604 71692
rect 179656 71680 179662 71732
rect 78674 71000 78680 71052
rect 78732 71040 78738 71052
rect 132034 71040 132040 71052
rect 78732 71012 132040 71040
rect 78732 71000 78738 71012
rect 132034 71000 132040 71012
rect 132092 71000 132098 71052
rect 138934 71000 138940 71052
rect 138992 71040 138998 71052
rect 152550 71040 152556 71052
rect 138992 71012 152556 71040
rect 138992 71000 138998 71012
rect 152550 71000 152556 71012
rect 152608 71000 152614 71052
rect 158346 71000 158352 71052
rect 158404 71040 158410 71052
rect 284386 71040 284392 71052
rect 158404 71012 284392 71040
rect 158404 71000 158410 71012
rect 284386 71000 284392 71012
rect 284444 71000 284450 71052
rect 138658 70320 138664 70372
rect 138716 70360 138722 70372
rect 142798 70360 142804 70372
rect 138716 70332 142804 70360
rect 138716 70320 138722 70332
rect 142798 70320 142804 70332
rect 142856 70320 142862 70372
rect 141510 70048 141516 70100
rect 141568 70088 141574 70100
rect 209866 70088 209872 70100
rect 141568 70060 209872 70088
rect 141568 70048 141574 70060
rect 209866 70048 209872 70060
rect 209924 70048 209930 70100
rect 155310 69980 155316 70032
rect 155368 70020 155374 70032
rect 382274 70020 382280 70032
rect 155368 69992 382280 70020
rect 155368 69980 155374 69992
rect 382274 69980 382280 69992
rect 382332 69980 382338 70032
rect 156598 69912 156604 69964
rect 156656 69952 156662 69964
rect 390554 69952 390560 69964
rect 156656 69924 390560 69952
rect 156656 69912 156662 69924
rect 390554 69912 390560 69924
rect 390612 69912 390618 69964
rect 171686 69844 171692 69896
rect 171744 69884 171750 69896
rect 426434 69884 426440 69896
rect 171744 69856 426440 69884
rect 171744 69844 171750 69856
rect 426434 69844 426440 69856
rect 426492 69844 426498 69896
rect 164878 69776 164884 69828
rect 164936 69816 164942 69828
rect 505094 69816 505100 69828
rect 164936 69788 505100 69816
rect 164936 69776 164942 69788
rect 505094 69776 505100 69788
rect 505152 69776 505158 69828
rect 166534 69708 166540 69760
rect 166592 69748 166598 69760
rect 518894 69748 518900 69760
rect 166592 69720 518900 69748
rect 166592 69708 166598 69720
rect 518894 69708 518900 69720
rect 518952 69708 518958 69760
rect 170306 69640 170312 69692
rect 170364 69680 170370 69692
rect 568574 69680 568580 69692
rect 170364 69652 568580 69680
rect 170364 69640 170370 69652
rect 568574 69640 568580 69652
rect 568632 69640 568638 69692
rect 170214 68960 170220 69012
rect 170272 69000 170278 69012
rect 171686 69000 171692 69012
rect 170272 68972 171692 69000
rect 170272 68960 170278 68972
rect 171686 68960 171692 68972
rect 171744 68960 171750 69012
rect 140038 68620 140044 68672
rect 140096 68660 140102 68672
rect 184934 68660 184940 68672
rect 140096 68632 184940 68660
rect 140096 68620 140102 68632
rect 184934 68620 184940 68632
rect 184992 68620 184998 68672
rect 142706 68552 142712 68604
rect 142764 68592 142770 68604
rect 218054 68592 218060 68604
rect 142764 68564 218060 68592
rect 142764 68552 142770 68564
rect 218054 68552 218060 68564
rect 218112 68552 218118 68604
rect 157058 68484 157064 68536
rect 157116 68524 157122 68536
rect 320174 68524 320180 68536
rect 157116 68496 320180 68524
rect 157116 68484 157122 68496
rect 320174 68484 320180 68496
rect 320232 68484 320238 68536
rect 153746 68416 153752 68468
rect 153804 68456 153810 68468
rect 362954 68456 362960 68468
rect 153804 68428 362960 68456
rect 153804 68416 153810 68428
rect 362954 68416 362960 68428
rect 363012 68416 363018 68468
rect 159266 68348 159272 68400
rect 159324 68388 159330 68400
rect 427814 68388 427820 68400
rect 159324 68360 427820 68388
rect 159324 68348 159330 68360
rect 427814 68348 427820 68360
rect 427872 68348 427878 68400
rect 169478 68280 169484 68332
rect 169536 68320 169542 68332
rect 564526 68320 564532 68332
rect 169536 68292 564532 68320
rect 169536 68280 169542 68292
rect 564526 68280 564532 68292
rect 564584 68280 564590 68332
rect 139946 67396 139952 67448
rect 140004 67436 140010 67448
rect 189074 67436 189080 67448
rect 140004 67408 189080 67436
rect 140004 67396 140010 67408
rect 189074 67396 189080 67408
rect 189132 67396 189138 67448
rect 147214 67328 147220 67380
rect 147272 67368 147278 67380
rect 270494 67368 270500 67380
rect 147272 67340 270500 67368
rect 147272 67328 147278 67340
rect 270494 67328 270500 67340
rect 270552 67328 270558 67380
rect 149698 67260 149704 67312
rect 149756 67300 149762 67312
rect 306374 67300 306380 67312
rect 149756 67272 306380 67300
rect 149756 67260 149762 67272
rect 306374 67260 306380 67272
rect 306432 67260 306438 67312
rect 160830 67192 160836 67244
rect 160888 67232 160894 67244
rect 347774 67232 347780 67244
rect 160888 67204 347780 67232
rect 160888 67192 160894 67204
rect 347774 67192 347780 67204
rect 347832 67192 347838 67244
rect 152458 67124 152464 67176
rect 152516 67164 152522 67176
rect 340966 67164 340972 67176
rect 152516 67136 340972 67164
rect 152516 67124 152522 67136
rect 340966 67124 340972 67136
rect 341024 67124 341030 67176
rect 159174 67056 159180 67108
rect 159232 67096 159238 67108
rect 437474 67096 437480 67108
rect 159232 67068 437480 67096
rect 159232 67056 159238 67068
rect 437474 67056 437480 67068
rect 437532 67056 437538 67108
rect 162026 66988 162032 67040
rect 162084 67028 162090 67040
rect 462314 67028 462320 67040
rect 162084 67000 462320 67028
rect 162084 66988 162090 67000
rect 462314 66988 462320 67000
rect 462372 66988 462378 67040
rect 167730 66920 167736 66972
rect 167788 66960 167794 66972
rect 539594 66960 539600 66972
rect 167788 66932 539600 66960
rect 167788 66920 167794 66932
rect 539594 66920 539600 66932
rect 539652 66920 539658 66972
rect 167638 66852 167644 66904
rect 167696 66892 167702 66904
rect 543734 66892 543740 66904
rect 167696 66864 543740 66892
rect 167696 66852 167702 66864
rect 543734 66852 543740 66864
rect 543792 66852 543798 66904
rect 137278 66172 137284 66224
rect 137336 66212 137342 66224
rect 140038 66212 140044 66224
rect 137336 66184 140044 66212
rect 137336 66172 137342 66184
rect 140038 66172 140044 66184
rect 140096 66172 140102 66224
rect 138566 66104 138572 66156
rect 138624 66144 138630 66156
rect 141510 66144 141516 66156
rect 138624 66116 141516 66144
rect 138624 66104 138630 66116
rect 141510 66104 141516 66116
rect 141568 66104 141574 66156
rect 141326 65900 141332 65952
rect 141384 65940 141390 65952
rect 202874 65940 202880 65952
rect 141384 65912 202880 65940
rect 141384 65900 141390 65912
rect 202874 65900 202880 65912
rect 202932 65900 202938 65952
rect 141418 65832 141424 65884
rect 141476 65872 141482 65884
rect 207014 65872 207020 65884
rect 141476 65844 207020 65872
rect 141476 65832 141482 65844
rect 207014 65832 207020 65844
rect 207072 65832 207078 65884
rect 142614 65764 142620 65816
rect 142672 65804 142678 65816
rect 220814 65804 220820 65816
rect 142672 65776 220820 65804
rect 142672 65764 142678 65776
rect 220814 65764 220820 65776
rect 220872 65764 220878 65816
rect 145466 65696 145472 65748
rect 145524 65736 145530 65748
rect 251266 65736 251272 65748
rect 145524 65708 251272 65736
rect 145524 65696 145530 65708
rect 251266 65696 251272 65708
rect 251324 65696 251330 65748
rect 145558 65628 145564 65680
rect 145616 65668 145622 65680
rect 256694 65668 256700 65680
rect 145616 65640 256700 65668
rect 145616 65628 145622 65640
rect 256694 65628 256700 65640
rect 256752 65628 256758 65680
rect 153654 65560 153660 65612
rect 153712 65600 153718 65612
rect 358814 65600 358820 65612
rect 153712 65572 358820 65600
rect 153712 65560 153718 65572
rect 358814 65560 358820 65572
rect 358872 65560 358878 65612
rect 102226 65492 102232 65544
rect 102284 65532 102290 65544
rect 125318 65532 125324 65544
rect 102284 65504 125324 65532
rect 102284 65492 102290 65504
rect 125318 65492 125324 65504
rect 125376 65492 125382 65544
rect 155218 65492 155224 65544
rect 155276 65532 155282 65544
rect 376754 65532 376760 65544
rect 155276 65504 376760 65532
rect 155276 65492 155282 65504
rect 376754 65492 376760 65504
rect 376812 65492 376818 65544
rect 144270 64472 144276 64524
rect 144328 64512 144334 64524
rect 234614 64512 234620 64524
rect 144328 64484 234620 64512
rect 144328 64472 144334 64484
rect 234614 64472 234620 64484
rect 234672 64472 234678 64524
rect 144178 64404 144184 64456
rect 144236 64444 144242 64456
rect 238754 64444 238760 64456
rect 144236 64416 238760 64444
rect 144236 64404 144242 64416
rect 238754 64404 238760 64416
rect 238812 64404 238818 64456
rect 148226 64336 148232 64388
rect 148284 64376 148290 64388
rect 292574 64376 292580 64388
rect 148284 64348 292580 64376
rect 148284 64336 148290 64348
rect 292574 64336 292580 64348
rect 292632 64336 292638 64388
rect 152366 64268 152372 64320
rect 152424 64308 152430 64320
rect 338114 64308 338120 64320
rect 152424 64280 338120 64308
rect 152424 64268 152430 64280
rect 338114 64268 338120 64280
rect 338172 64268 338178 64320
rect 162578 64200 162584 64252
rect 162636 64240 162642 64252
rect 368474 64240 368480 64252
rect 162636 64212 368480 64240
rect 162636 64200 162642 64212
rect 368474 64200 368480 64212
rect 368532 64200 368538 64252
rect 169018 64132 169024 64184
rect 169076 64172 169082 64184
rect 561674 64172 561680 64184
rect 169076 64144 561680 64172
rect 169076 64132 169082 64144
rect 561674 64132 561680 64144
rect 561732 64132 561738 64184
rect 147030 63112 147036 63164
rect 147088 63152 147094 63164
rect 274634 63152 274640 63164
rect 147088 63124 274640 63152
rect 147088 63112 147094 63124
rect 274634 63112 274640 63124
rect 274692 63112 274698 63164
rect 149606 63044 149612 63096
rect 149664 63084 149670 63096
rect 309134 63084 309140 63096
rect 149664 63056 309140 63084
rect 149664 63044 149670 63056
rect 309134 63044 309140 63056
rect 309192 63044 309198 63096
rect 155126 62976 155132 63028
rect 155184 63016 155190 63028
rect 373994 63016 374000 63028
rect 155184 62988 374000 63016
rect 155184 62976 155190 62988
rect 373994 62976 374000 62988
rect 374052 62976 374058 63028
rect 157978 62908 157984 62960
rect 158036 62948 158042 62960
rect 408494 62948 408500 62960
rect 158036 62920 408500 62948
rect 158036 62908 158042 62920
rect 408494 62908 408500 62920
rect 408552 62908 408558 62960
rect 163590 62840 163596 62892
rect 163648 62880 163654 62892
rect 488534 62880 488540 62892
rect 163648 62852 488540 62880
rect 163648 62840 163654 62852
rect 488534 62840 488540 62852
rect 488592 62840 488598 62892
rect 168926 62772 168932 62824
rect 168984 62812 168990 62824
rect 557534 62812 557540 62824
rect 168984 62784 557540 62812
rect 168984 62772 168990 62784
rect 557534 62772 557540 62784
rect 557592 62772 557598 62824
rect 139854 61480 139860 61532
rect 139912 61520 139918 61532
rect 185026 61520 185032 61532
rect 139912 61492 185032 61520
rect 139912 61480 139918 61492
rect 185026 61480 185032 61492
rect 185084 61480 185090 61532
rect 157886 61412 157892 61464
rect 157944 61452 157950 61464
rect 412634 61452 412640 61464
rect 157944 61424 412640 61452
rect 157944 61412 157950 61424
rect 412634 61412 412640 61424
rect 412692 61412 412698 61464
rect 166350 61344 166356 61396
rect 166408 61384 166414 61396
rect 525794 61384 525800 61396
rect 166408 61356 525800 61384
rect 166408 61344 166414 61356
rect 525794 61344 525800 61356
rect 525852 61344 525858 61396
rect 118510 60664 118516 60716
rect 118568 60704 118574 60716
rect 580166 60704 580172 60716
rect 118568 60676 580172 60704
rect 118568 60664 118574 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 137186 59984 137192 60036
rect 137244 60024 137250 60036
rect 138658 60024 138664 60036
rect 137244 59996 138664 60024
rect 137244 59984 137250 59996
rect 138658 59984 138664 59996
rect 138716 59984 138722 60036
rect 159082 59984 159088 60036
rect 159140 60024 159146 60036
rect 433334 60024 433340 60036
rect 159140 59996 433340 60024
rect 159140 59984 159146 59996
rect 433334 59984 433340 59996
rect 433392 59984 433398 60036
rect 156506 58624 156512 58676
rect 156564 58664 156570 58676
rect 401594 58664 401600 58676
rect 156564 58636 401600 58664
rect 156564 58624 156570 58636
rect 401594 58624 401600 58636
rect 401652 58624 401658 58676
rect 163498 57264 163504 57316
rect 163556 57304 163562 57316
rect 481634 57304 481640 57316
rect 163556 57276 481640 57304
rect 163556 57264 163562 57276
rect 481634 57264 481640 57276
rect 481692 57264 481698 57316
rect 164786 57196 164792 57248
rect 164844 57236 164850 57248
rect 507854 57236 507860 57248
rect 164844 57208 507860 57236
rect 164844 57196 164850 57208
rect 507854 57196 507860 57208
rect 507912 57196 507918 57248
rect 95234 53048 95240 53100
rect 95292 53088 95298 53100
rect 125226 53088 125232 53100
rect 95292 53060 125232 53088
rect 95292 53048 95298 53060
rect 125226 53048 125232 53060
rect 125284 53048 125290 53100
rect 182818 46860 182824 46912
rect 182876 46900 182882 46912
rect 580166 46900 580172 46912
rect 182876 46872 580172 46900
rect 182876 46860 182882 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 139762 46180 139768 46232
rect 139820 46220 139826 46232
rect 180794 46220 180800 46232
rect 139820 46192 180800 46220
rect 139820 46180 139826 46192
rect 180794 46180 180800 46192
rect 180852 46180 180858 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 174078 45540 174084 45552
rect 3476 45512 174084 45540
rect 3476 45500 3482 45512
rect 174078 45500 174084 45512
rect 174136 45500 174142 45552
rect 135990 44956 135996 45008
rect 136048 44996 136054 45008
rect 142614 44996 142620 45008
rect 136048 44968 142620 44996
rect 136048 44956 136054 44968
rect 142614 44956 142620 44968
rect 142672 44956 142678 45008
rect 70394 44888 70400 44940
rect 70452 44928 70458 44940
rect 130286 44928 130292 44940
rect 70452 44900 130292 44928
rect 70452 44888 70458 44900
rect 130286 44888 130292 44900
rect 130344 44888 130350 44940
rect 34514 44820 34520 44872
rect 34572 44860 34578 44872
rect 127342 44860 127348 44872
rect 34572 44832 127348 44860
rect 34572 44820 34578 44832
rect 127342 44820 127348 44832
rect 127400 44820 127406 44872
rect 138474 44820 138480 44872
rect 138532 44860 138538 44872
rect 147030 44860 147036 44872
rect 138532 44832 147036 44860
rect 138532 44820 138538 44832
rect 147030 44820 147036 44832
rect 147088 44820 147094 44872
rect 171594 43392 171600 43444
rect 171652 43432 171658 43444
rect 411254 43432 411260 43444
rect 171652 43404 411260 43432
rect 171652 43392 171658 43404
rect 411254 43392 411260 43404
rect 411312 43392 411318 43444
rect 19334 42032 19340 42084
rect 19392 42072 19398 42084
rect 125134 42072 125140 42084
rect 19392 42044 125140 42072
rect 19392 42032 19398 42044
rect 125134 42032 125140 42044
rect 125192 42032 125198 42084
rect 162210 42032 162216 42084
rect 162268 42072 162274 42084
rect 390646 42072 390652 42084
rect 162268 42044 390652 42072
rect 162268 42032 162274 42044
rect 390646 42032 390652 42044
rect 390704 42032 390710 42084
rect 172422 40672 172428 40724
rect 172480 40712 172486 40724
rect 418154 40712 418160 40724
rect 172480 40684 418160 40712
rect 172480 40672 172486 40684
rect 418154 40672 418160 40684
rect 418212 40672 418218 40724
rect 120074 40264 120080 40316
rect 120132 40304 120138 40316
rect 123478 40304 123484 40316
rect 120132 40276 123484 40304
rect 120132 40264 120138 40276
rect 123478 40264 123484 40276
rect 123536 40264 123542 40316
rect 172330 39312 172336 39364
rect 172388 39352 172394 39364
rect 404354 39352 404360 39364
rect 172388 39324 404360 39352
rect 172388 39312 172394 39324
rect 404354 39312 404360 39324
rect 404412 39312 404418 39364
rect 172238 37884 172244 37936
rect 172296 37924 172302 37936
rect 397454 37924 397460 37936
rect 172296 37896 397460 37924
rect 172296 37884 172302 37896
rect 397454 37884 397460 37896
rect 397512 37884 397518 37936
rect 88334 36524 88340 36576
rect 88392 36564 88398 36576
rect 125042 36564 125048 36576
rect 88392 36536 125048 36564
rect 88392 36524 88398 36536
rect 125042 36524 125048 36536
rect 125100 36524 125106 36576
rect 145374 35572 145380 35624
rect 145432 35612 145438 35624
rect 259454 35612 259460 35624
rect 145432 35584 259460 35612
rect 145432 35572 145438 35584
rect 259454 35572 259460 35584
rect 259512 35572 259518 35624
rect 146938 35504 146944 35556
rect 146996 35544 147002 35556
rect 276014 35544 276020 35556
rect 146996 35516 276020 35544
rect 146996 35504 147002 35516
rect 276014 35504 276020 35516
rect 276072 35504 276078 35556
rect 148134 35436 148140 35488
rect 148192 35476 148198 35488
rect 287054 35476 287060 35488
rect 148192 35448 287060 35476
rect 148192 35436 148198 35448
rect 287054 35436 287060 35448
rect 287112 35436 287118 35488
rect 148042 35368 148048 35420
rect 148100 35408 148106 35420
rect 293954 35408 293960 35420
rect 148100 35380 293960 35408
rect 148100 35368 148106 35380
rect 293954 35368 293960 35380
rect 294012 35368 294018 35420
rect 149514 35300 149520 35352
rect 149572 35340 149578 35352
rect 304994 35340 305000 35352
rect 149572 35312 305000 35340
rect 149572 35300 149578 35312
rect 304994 35300 305000 35312
rect 305052 35300 305058 35352
rect 149422 35232 149428 35284
rect 149480 35272 149486 35284
rect 307754 35272 307760 35284
rect 149480 35244 307760 35272
rect 149480 35232 149486 35244
rect 307754 35232 307760 35244
rect 307812 35232 307818 35284
rect 159726 35164 159732 35216
rect 159784 35204 159790 35216
rect 382366 35204 382372 35216
rect 159784 35176 382372 35204
rect 159784 35164 159790 35176
rect 382366 35164 382372 35176
rect 382424 35164 382430 35216
rect 139670 34076 139676 34128
rect 139728 34116 139734 34128
rect 187694 34116 187700 34128
rect 139728 34088 187700 34116
rect 139728 34076 139734 34088
rect 187694 34076 187700 34088
rect 187752 34076 187758 34128
rect 141142 34008 141148 34060
rect 141200 34048 141206 34060
rect 198734 34048 198740 34060
rect 141200 34020 198740 34048
rect 141200 34008 141206 34020
rect 198734 34008 198740 34020
rect 198792 34008 198798 34060
rect 141050 33940 141056 33992
rect 141108 33980 141114 33992
rect 201494 33980 201500 33992
rect 141108 33952 201500 33980
rect 141108 33940 141114 33952
rect 201494 33940 201500 33952
rect 201552 33940 201558 33992
rect 141234 33872 141240 33924
rect 141292 33912 141298 33924
rect 205634 33912 205640 33924
rect 141292 33884 205640 33912
rect 141292 33872 141298 33884
rect 205634 33872 205640 33884
rect 205692 33872 205698 33924
rect 144086 33804 144092 33856
rect 144144 33844 144150 33856
rect 234706 33844 234712 33856
rect 144144 33816 234712 33844
rect 144144 33804 144150 33816
rect 234706 33804 234712 33816
rect 234764 33804 234770 33856
rect 146846 33736 146852 33788
rect 146904 33776 146910 33788
rect 269114 33776 269120 33788
rect 146904 33748 269120 33776
rect 146904 33736 146910 33748
rect 269114 33736 269120 33748
rect 269172 33736 269178 33788
rect 171686 33056 171692 33108
rect 171744 33096 171750 33108
rect 580166 33096 580172 33108
rect 171744 33068 580172 33096
rect 171744 33056 171750 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 180886 33028 180892 33040
rect 3476 33000 180892 33028
rect 3476 32988 3482 33000
rect 180886 32988 180892 33000
rect 180944 32988 180950 33040
rect 156414 32716 156420 32768
rect 156472 32756 156478 32768
rect 391934 32756 391940 32768
rect 156472 32728 391940 32756
rect 156472 32716 156478 32728
rect 391934 32716 391940 32728
rect 391992 32716 391998 32768
rect 160002 32648 160008 32700
rect 160060 32688 160066 32700
rect 434714 32688 434720 32700
rect 160060 32660 434720 32688
rect 160060 32648 160066 32660
rect 434714 32648 434720 32660
rect 434772 32648 434778 32700
rect 161934 32580 161940 32632
rect 161992 32620 161998 32632
rect 463694 32620 463700 32632
rect 161992 32592 463700 32620
rect 161992 32580 161998 32592
rect 463694 32580 463700 32592
rect 463752 32580 463758 32632
rect 163406 32512 163412 32564
rect 163464 32552 163470 32564
rect 481726 32552 481732 32564
rect 163464 32524 481732 32552
rect 163464 32512 163470 32524
rect 481726 32512 481732 32524
rect 481784 32512 481790 32564
rect 167546 32444 167552 32496
rect 167604 32484 167610 32496
rect 539686 32484 539692 32496
rect 167604 32456 539692 32484
rect 167604 32444 167610 32456
rect 539686 32444 539692 32456
rect 539744 32444 539750 32496
rect 170122 32376 170128 32428
rect 170180 32416 170186 32428
rect 574094 32416 574100 32428
rect 170180 32388 574100 32416
rect 170180 32376 170186 32388
rect 574094 32376 574100 32388
rect 574152 32376 574158 32428
rect 143994 31424 144000 31476
rect 144052 31464 144058 31476
rect 242894 31464 242900 31476
rect 144052 31436 242900 31464
rect 144052 31424 144058 31436
rect 242894 31424 242900 31436
rect 242952 31424 242958 31476
rect 146754 31356 146760 31408
rect 146812 31396 146818 31408
rect 267826 31396 267832 31408
rect 146812 31368 267832 31396
rect 146812 31356 146818 31368
rect 267826 31356 267832 31368
rect 267884 31356 267890 31408
rect 147950 31288 147956 31340
rect 148008 31328 148014 31340
rect 289814 31328 289820 31340
rect 148008 31300 289820 31328
rect 148008 31288 148014 31300
rect 289814 31288 289820 31300
rect 289872 31288 289878 31340
rect 154114 31220 154120 31272
rect 154172 31260 154178 31272
rect 332594 31260 332600 31272
rect 154172 31232 332600 31260
rect 154172 31220 154178 31232
rect 332594 31220 332600 31232
rect 332652 31220 332658 31272
rect 153562 31152 153568 31204
rect 153620 31192 153626 31204
rect 357526 31192 357532 31204
rect 153620 31164 357532 31192
rect 153620 31152 153626 31164
rect 357526 31152 357532 31164
rect 357584 31152 357590 31204
rect 156966 31084 156972 31136
rect 157024 31124 157030 31136
rect 389174 31124 389180 31136
rect 157024 31096 389180 31124
rect 157024 31084 157030 31096
rect 389174 31084 389180 31096
rect 389232 31084 389238 31136
rect 166258 31016 166264 31068
rect 166316 31056 166322 31068
rect 524414 31056 524420 31068
rect 166316 31028 524420 31056
rect 166316 31016 166322 31028
rect 524414 31016 524420 31028
rect 524472 31016 524478 31068
rect 140866 30064 140872 30116
rect 140924 30104 140930 30116
rect 204254 30104 204260 30116
rect 140924 30076 204260 30104
rect 140924 30064 140930 30076
rect 204254 30064 204260 30076
rect 204312 30064 204318 30116
rect 140958 29996 140964 30048
rect 141016 30036 141022 30048
rect 208394 30036 208400 30048
rect 141016 30008 208400 30036
rect 141016 29996 141022 30008
rect 208394 29996 208400 30008
rect 208452 29996 208458 30048
rect 143902 29928 143908 29980
rect 143960 29968 143966 29980
rect 233234 29968 233240 29980
rect 143960 29940 233240 29968
rect 143960 29928 143966 29940
rect 233234 29928 233240 29940
rect 233292 29928 233298 29980
rect 143810 29860 143816 29912
rect 143868 29900 143874 29912
rect 235994 29900 236000 29912
rect 143868 29872 236000 29900
rect 143868 29860 143874 29872
rect 235994 29860 236000 29872
rect 236052 29860 236058 29912
rect 145282 29792 145288 29844
rect 145340 29832 145346 29844
rect 253934 29832 253940 29844
rect 145340 29804 253940 29832
rect 145340 29792 145346 29804
rect 253934 29792 253940 29804
rect 253992 29792 253998 29844
rect 145190 29724 145196 29776
rect 145248 29764 145254 29776
rect 258074 29764 258080 29776
rect 145248 29736 258080 29764
rect 145248 29724 145254 29736
rect 258074 29724 258080 29736
rect 258132 29724 258138 29776
rect 166166 29656 166172 29708
rect 166224 29696 166230 29708
rect 521654 29696 521660 29708
rect 166224 29668 521660 29696
rect 166224 29656 166230 29668
rect 521654 29656 521660 29668
rect 521712 29656 521718 29708
rect 167454 29588 167460 29640
rect 167512 29628 167518 29640
rect 542354 29628 542360 29640
rect 167512 29600 542360 29628
rect 167512 29588 167518 29600
rect 542354 29588 542360 29600
rect 542412 29588 542418 29640
rect 148686 28500 148692 28552
rect 148744 28540 148750 28552
rect 190454 28540 190460 28552
rect 148744 28512 190460 28540
rect 148744 28500 148750 28512
rect 190454 28500 190460 28512
rect 190512 28500 190518 28552
rect 139578 28432 139584 28484
rect 139636 28472 139642 28484
rect 186314 28472 186320 28484
rect 139636 28444 186320 28472
rect 139636 28432 139642 28444
rect 186314 28432 186320 28444
rect 186372 28432 186378 28484
rect 140774 28364 140780 28416
rect 140832 28404 140838 28416
rect 201586 28404 201592 28416
rect 140832 28376 201592 28404
rect 140832 28364 140838 28376
rect 201586 28364 201592 28376
rect 201644 28364 201650 28416
rect 146662 28296 146668 28348
rect 146720 28336 146726 28348
rect 271874 28336 271880 28348
rect 146720 28308 271880 28336
rect 146720 28296 146726 28308
rect 271874 28296 271880 28308
rect 271932 28296 271938 28348
rect 147858 28228 147864 28280
rect 147916 28268 147922 28280
rect 285674 28268 285680 28280
rect 147916 28240 285680 28268
rect 147916 28228 147922 28240
rect 285674 28228 285680 28240
rect 285732 28228 285738 28280
rect 322198 28228 322204 28280
rect 322256 28268 322262 28280
rect 580994 28268 581000 28280
rect 322256 28240 581000 28268
rect 322256 28228 322262 28240
rect 580994 28228 581000 28240
rect 581052 28228 581058 28280
rect 140498 27276 140504 27328
rect 140556 27316 140562 27328
rect 176746 27316 176752 27328
rect 140556 27288 176752 27316
rect 140556 27276 140562 27288
rect 176746 27276 176752 27288
rect 176804 27276 176810 27328
rect 139394 27208 139400 27260
rect 139452 27248 139458 27260
rect 179414 27248 179420 27260
rect 139452 27220 179420 27248
rect 139452 27208 139458 27220
rect 179414 27208 179420 27220
rect 179472 27208 179478 27260
rect 139486 27140 139492 27192
rect 139544 27180 139550 27192
rect 183554 27180 183560 27192
rect 139544 27152 183560 27180
rect 139544 27140 139550 27152
rect 183554 27140 183560 27152
rect 183612 27140 183618 27192
rect 146570 27072 146576 27124
rect 146628 27112 146634 27124
rect 276106 27112 276112 27124
rect 146628 27084 276112 27112
rect 146628 27072 146634 27084
rect 276106 27072 276112 27084
rect 276164 27072 276170 27124
rect 149330 27004 149336 27056
rect 149388 27044 149394 27056
rect 310514 27044 310520 27056
rect 149388 27016 310520 27044
rect 149388 27004 149394 27016
rect 310514 27004 310520 27016
rect 310572 27004 310578 27056
rect 152274 26936 152280 26988
rect 152332 26976 152338 26988
rect 339494 26976 339500 26988
rect 152332 26948 339500 26976
rect 152332 26936 152338 26948
rect 339494 26936 339500 26948
rect 339552 26936 339558 26988
rect 164694 26868 164700 26920
rect 164752 26908 164758 26920
rect 506474 26908 506480 26920
rect 164752 26880 506480 26908
rect 164752 26868 164758 26880
rect 506474 26868 506480 26880
rect 506532 26868 506538 26920
rect 142522 25984 142528 26036
rect 142580 26024 142586 26036
rect 222194 26024 222200 26036
rect 142580 25996 222200 26024
rect 142580 25984 142586 25996
rect 222194 25984 222200 25996
rect 222252 25984 222258 26036
rect 146478 25916 146484 25968
rect 146536 25956 146542 25968
rect 278774 25956 278780 25968
rect 146536 25928 278780 25956
rect 146536 25916 146542 25928
rect 278774 25916 278780 25928
rect 278832 25916 278838 25968
rect 149238 25848 149244 25900
rect 149296 25888 149302 25900
rect 307846 25888 307852 25900
rect 149296 25860 307852 25888
rect 149296 25848 149302 25860
rect 307846 25848 307852 25860
rect 307904 25848 307910 25900
rect 152182 25780 152188 25832
rect 152240 25820 152246 25832
rect 346394 25820 346400 25832
rect 152240 25792 346400 25820
rect 152240 25780 152246 25792
rect 346394 25780 346400 25792
rect 346452 25780 346458 25832
rect 166074 25712 166080 25764
rect 166132 25752 166138 25764
rect 517514 25752 517520 25764
rect 166132 25724 517520 25752
rect 166132 25712 166138 25724
rect 517514 25712 517520 25724
rect 517572 25712 517578 25764
rect 170674 25644 170680 25696
rect 170732 25684 170738 25696
rect 558914 25684 558920 25696
rect 170732 25656 558920 25684
rect 170732 25644 170738 25656
rect 558914 25644 558920 25656
rect 558972 25644 558978 25696
rect 168834 25576 168840 25628
rect 168892 25616 168898 25628
rect 563054 25616 563060 25628
rect 168892 25588 563060 25616
rect 168892 25576 168898 25588
rect 563054 25576 563060 25588
rect 563112 25576 563118 25628
rect 170030 25508 170036 25560
rect 170088 25548 170094 25560
rect 572714 25548 572720 25560
rect 170088 25520 572720 25548
rect 170088 25508 170094 25520
rect 572714 25508 572720 25520
rect 572772 25508 572778 25560
rect 142338 24556 142344 24608
rect 142396 24596 142402 24608
rect 215294 24596 215300 24608
rect 142396 24568 215300 24596
rect 142396 24556 142402 24568
rect 215294 24556 215300 24568
rect 215352 24556 215358 24608
rect 142430 24488 142436 24540
rect 142488 24528 142494 24540
rect 218146 24528 218152 24540
rect 142488 24500 218152 24528
rect 142488 24488 142494 24500
rect 218146 24488 218152 24500
rect 218204 24488 218210 24540
rect 147766 24420 147772 24472
rect 147824 24460 147830 24472
rect 292666 24460 292672 24472
rect 147824 24432 292672 24460
rect 147824 24420 147830 24432
rect 292666 24420 292672 24432
rect 292724 24420 292730 24472
rect 155034 24352 155040 24404
rect 155092 24392 155098 24404
rect 374086 24392 374092 24404
rect 155092 24364 374092 24392
rect 155092 24352 155098 24364
rect 374086 24352 374092 24364
rect 374144 24352 374150 24404
rect 167362 24284 167368 24336
rect 167420 24324 167426 24336
rect 467098 24324 467104 24336
rect 167420 24296 467104 24324
rect 167420 24284 167426 24296
rect 467098 24284 467104 24296
rect 467156 24284 467162 24336
rect 167270 24216 167276 24268
rect 167328 24256 167334 24268
rect 535454 24256 535460 24268
rect 167328 24228 535460 24256
rect 167328 24216 167334 24228
rect 535454 24216 535460 24228
rect 535512 24216 535518 24268
rect 167178 24148 167184 24200
rect 167236 24188 167242 24200
rect 538214 24188 538220 24200
rect 167236 24160 538220 24188
rect 167236 24148 167242 24160
rect 538214 24148 538220 24160
rect 538272 24148 538278 24200
rect 168742 24080 168748 24132
rect 168800 24120 168806 24132
rect 552014 24120 552020 24132
rect 168800 24092 552020 24120
rect 168800 24080 168806 24092
rect 552014 24080 552020 24092
rect 552072 24080 552078 24132
rect 149146 23332 149152 23384
rect 149204 23372 149210 23384
rect 303614 23372 303620 23384
rect 149204 23344 303620 23372
rect 149204 23332 149210 23344
rect 303614 23332 303620 23344
rect 303672 23332 303678 23384
rect 3418 23264 3424 23316
rect 3476 23304 3482 23316
rect 173986 23304 173992 23316
rect 3476 23276 173992 23304
rect 3476 23264 3482 23276
rect 173986 23264 173992 23276
rect 174044 23264 174050 23316
rect 153470 23196 153476 23248
rect 153528 23236 153534 23248
rect 360194 23236 360200 23248
rect 153528 23208 360200 23236
rect 153528 23196 153534 23208
rect 360194 23196 360200 23208
rect 360252 23196 360258 23248
rect 154942 23128 154948 23180
rect 155000 23168 155006 23180
rect 379514 23168 379520 23180
rect 155000 23140 379520 23168
rect 155000 23128 155006 23140
rect 379514 23128 379520 23140
rect 379572 23128 379578 23180
rect 164510 23060 164516 23112
rect 164568 23100 164574 23112
rect 498286 23100 498292 23112
rect 164568 23072 498292 23100
rect 164568 23060 164574 23072
rect 498286 23060 498292 23072
rect 498344 23060 498350 23112
rect 164602 22992 164608 23044
rect 164660 23032 164666 23044
rect 509234 23032 509240 23044
rect 164660 23004 509240 23032
rect 164660 22992 164666 23004
rect 509234 22992 509240 23004
rect 509292 22992 509298 23044
rect 165890 22924 165896 22976
rect 165948 22964 165954 22976
rect 516134 22964 516140 22976
rect 165948 22936 516140 22964
rect 165948 22924 165954 22936
rect 516134 22924 516140 22936
rect 516192 22924 516198 22976
rect 165982 22856 165988 22908
rect 166040 22896 166046 22908
rect 520274 22896 520280 22908
rect 166040 22868 520280 22896
rect 166040 22856 166046 22868
rect 520274 22856 520280 22868
rect 520332 22856 520338 22908
rect 74534 22788 74540 22840
rect 74592 22828 74598 22840
rect 128446 22828 128452 22840
rect 74592 22800 128452 22828
rect 74592 22788 74598 22800
rect 128446 22788 128452 22800
rect 128504 22788 128510 22840
rect 168650 22788 168656 22840
rect 168708 22828 168714 22840
rect 556154 22828 556160 22840
rect 168708 22800 556160 22828
rect 168708 22788 168714 22800
rect 556154 22788 556160 22800
rect 556212 22788 556218 22840
rect 118418 22720 118424 22772
rect 118476 22760 118482 22772
rect 580166 22760 580172 22772
rect 118476 22732 580172 22760
rect 118476 22720 118482 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 152090 21632 152096 21684
rect 152148 21672 152154 21684
rect 343634 21672 343640 21684
rect 152148 21644 343640 21672
rect 152148 21632 152154 21644
rect 343634 21632 343640 21644
rect 343692 21632 343698 21684
rect 160646 21564 160652 21616
rect 160704 21604 160710 21616
rect 447134 21604 447140 21616
rect 160704 21576 447140 21604
rect 160704 21564 160710 21576
rect 447134 21564 447140 21576
rect 447192 21564 447198 21616
rect 161842 21496 161848 21548
rect 161900 21536 161906 21548
rect 473354 21536 473360 21548
rect 161900 21508 473360 21536
rect 161900 21496 161906 21508
rect 473354 21496 473360 21508
rect 473412 21496 473418 21548
rect 163314 21428 163320 21480
rect 163372 21468 163378 21480
rect 484394 21468 484400 21480
rect 163372 21440 484400 21468
rect 163372 21428 163378 21440
rect 484394 21428 484400 21440
rect 484452 21428 484458 21480
rect 124306 21360 124312 21412
rect 124364 21400 124370 21412
rect 134334 21400 134340 21412
rect 124364 21372 134340 21400
rect 124364 21360 124370 21372
rect 134334 21360 134340 21372
rect 134392 21360 134398 21412
rect 164418 21360 164424 21412
rect 164476 21400 164482 21412
rect 506566 21400 506572 21412
rect 164476 21372 506572 21400
rect 164476 21360 164482 21372
rect 506566 21360 506572 21372
rect 506624 21360 506630 21412
rect 145006 20340 145012 20392
rect 145064 20380 145070 20392
rect 255314 20380 255320 20392
rect 145064 20352 255320 20380
rect 145064 20340 145070 20352
rect 255314 20340 255320 20352
rect 255372 20340 255378 20392
rect 145098 20272 145104 20324
rect 145156 20312 145162 20324
rect 262214 20312 262220 20324
rect 145156 20284 262220 20312
rect 145156 20272 145162 20284
rect 262214 20272 262220 20284
rect 262272 20272 262278 20324
rect 146386 20204 146392 20256
rect 146444 20244 146450 20256
rect 273254 20244 273260 20256
rect 146444 20216 273260 20244
rect 146444 20204 146450 20216
rect 273254 20204 273260 20216
rect 273312 20204 273318 20256
rect 247678 20136 247684 20188
rect 247736 20176 247742 20188
rect 456794 20176 456800 20188
rect 247736 20148 456800 20176
rect 247736 20136 247742 20148
rect 456794 20136 456800 20148
rect 456852 20136 456858 20188
rect 138382 20068 138388 20120
rect 138440 20108 138446 20120
rect 162854 20108 162860 20120
rect 138440 20080 162860 20108
rect 138440 20068 138446 20080
rect 162854 20068 162860 20080
rect 162912 20068 162918 20120
rect 253198 20068 253204 20120
rect 253256 20108 253262 20120
rect 465074 20108 465080 20120
rect 253256 20080 465080 20108
rect 253256 20068 253262 20080
rect 465074 20068 465080 20080
rect 465132 20068 465138 20120
rect 85574 20000 85580 20052
rect 85632 20040 85638 20052
rect 131666 20040 131672 20052
rect 85632 20012 131672 20040
rect 85632 20000 85638 20012
rect 131666 20000 131672 20012
rect 131724 20000 131730 20052
rect 160554 20000 160560 20052
rect 160612 20040 160618 20052
rect 455414 20040 455420 20052
rect 160612 20012 455420 20040
rect 160612 20000 160618 20012
rect 455414 20000 455420 20012
rect 455472 20000 455478 20052
rect 45554 19932 45560 19984
rect 45612 19972 45618 19984
rect 120810 19972 120816 19984
rect 45612 19944 120816 19972
rect 45612 19932 45618 19944
rect 120810 19932 120816 19944
rect 120868 19932 120874 19984
rect 161750 19932 161756 19984
rect 161808 19972 161814 19984
rect 465166 19972 465172 19984
rect 161808 19944 465172 19972
rect 161808 19932 161814 19944
rect 465166 19932 465172 19944
rect 465224 19932 465230 19984
rect 160462 18844 160468 18896
rect 160520 18884 160526 18896
rect 448514 18884 448520 18896
rect 160520 18856 448520 18884
rect 160520 18844 160526 18856
rect 448514 18844 448520 18856
rect 448572 18844 448578 18896
rect 160370 18776 160376 18828
rect 160428 18816 160434 18828
rect 451274 18816 451280 18828
rect 160428 18788 451280 18816
rect 160428 18776 160434 18788
rect 451274 18776 451280 18788
rect 451332 18776 451338 18828
rect 117314 18708 117320 18760
rect 117372 18748 117378 18760
rect 134242 18748 134248 18760
rect 117372 18720 134248 18748
rect 117372 18708 117378 18720
rect 134242 18708 134248 18720
rect 134300 18708 134306 18760
rect 168466 18708 168472 18760
rect 168524 18748 168530 18760
rect 553394 18748 553400 18760
rect 168524 18720 553400 18748
rect 168524 18708 168530 18720
rect 553394 18708 553400 18720
rect 553452 18708 553458 18760
rect 31754 18640 31760 18692
rect 31812 18680 31818 18692
rect 122282 18680 122288 18692
rect 31812 18652 122288 18680
rect 31812 18640 31818 18652
rect 122282 18640 122288 18652
rect 122340 18640 122346 18692
rect 168374 18640 168380 18692
rect 168432 18680 168438 18692
rect 556246 18680 556252 18692
rect 168432 18652 556252 18680
rect 168432 18640 168438 18652
rect 556246 18640 556252 18652
rect 556304 18640 556310 18692
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 126238 18612 126244 18624
rect 4212 18584 126244 18612
rect 4212 18572 4218 18584
rect 126238 18572 126244 18584
rect 126296 18572 126302 18624
rect 168558 18572 168564 18624
rect 168616 18612 168622 18624
rect 560294 18612 560300 18624
rect 168616 18584 560300 18612
rect 168616 18572 168622 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 157702 17552 157708 17604
rect 157760 17592 157766 17604
rect 415394 17592 415400 17604
rect 157760 17564 415400 17592
rect 157760 17552 157766 17564
rect 415394 17552 415400 17564
rect 415452 17552 415458 17604
rect 157794 17484 157800 17536
rect 157852 17524 157858 17536
rect 419534 17524 419540 17536
rect 157852 17496 419540 17524
rect 157852 17484 157858 17496
rect 419534 17484 419540 17496
rect 419592 17484 419598 17536
rect 171962 17416 171968 17468
rect 172020 17456 172026 17468
rect 440234 17456 440240 17468
rect 172020 17428 440240 17456
rect 172020 17416 172026 17428
rect 440234 17416 440240 17428
rect 440292 17416 440298 17468
rect 160278 17348 160284 17400
rect 160336 17388 160342 17400
rect 448606 17388 448612 17400
rect 160336 17360 448612 17388
rect 160336 17348 160342 17360
rect 448606 17348 448612 17360
rect 448664 17348 448670 17400
rect 163222 17280 163228 17332
rect 163280 17320 163286 17332
rect 492674 17320 492680 17332
rect 163280 17292 492680 17320
rect 163280 17280 163286 17292
rect 492674 17280 492680 17292
rect 492732 17280 492738 17332
rect 167086 17212 167092 17264
rect 167144 17252 167150 17264
rect 545114 17252 545120 17264
rect 167144 17224 545120 17252
rect 167144 17212 167150 17224
rect 545114 17212 545120 17224
rect 545172 17212 545178 17264
rect 154850 16124 154856 16176
rect 154908 16164 154914 16176
rect 378410 16164 378416 16176
rect 154908 16136 378416 16164
rect 154908 16124 154914 16136
rect 378410 16124 378416 16136
rect 378468 16124 378474 16176
rect 156322 16056 156328 16108
rect 156380 16096 156386 16108
rect 395338 16096 395344 16108
rect 156380 16068 395344 16096
rect 156380 16056 156386 16068
rect 395338 16056 395344 16068
rect 395396 16056 395402 16108
rect 156230 15988 156236 16040
rect 156288 16028 156294 16040
rect 398834 16028 398840 16040
rect 156288 16000 398840 16028
rect 156288 15988 156294 16000
rect 398834 15988 398840 16000
rect 398892 15988 398898 16040
rect 174538 15920 174544 15972
rect 174596 15960 174602 15972
rect 425698 15960 425704 15972
rect 174596 15932 425704 15960
rect 174596 15920 174602 15932
rect 425698 15920 425704 15932
rect 425756 15920 425762 15972
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 124950 15892 124956 15904
rect 14332 15864 124956 15892
rect 14332 15852 14338 15864
rect 124950 15852 124956 15864
rect 125008 15852 125014 15904
rect 167914 15852 167920 15904
rect 167972 15892 167978 15904
rect 541986 15892 541992 15904
rect 167972 15864 541992 15892
rect 167972 15852 167978 15864
rect 541986 15852 541992 15864
rect 542044 15852 542050 15904
rect 143718 14764 143724 14816
rect 143776 14804 143782 14816
rect 241698 14804 241704 14816
rect 143776 14776 241704 14804
rect 143776 14764 143782 14776
rect 241698 14764 241704 14776
rect 241756 14764 241762 14816
rect 154666 14696 154672 14748
rect 154724 14736 154730 14748
rect 381170 14736 381176 14748
rect 154724 14708 381176 14736
rect 154724 14696 154730 14708
rect 381170 14696 381176 14708
rect 381228 14696 381234 14748
rect 154758 14628 154764 14680
rect 154816 14668 154822 14680
rect 384298 14668 384304 14680
rect 154816 14640 384304 14668
rect 154816 14628 154822 14640
rect 384298 14628 384304 14640
rect 384356 14628 384362 14680
rect 154574 14560 154580 14612
rect 154632 14600 154638 14612
rect 385954 14600 385960 14612
rect 154632 14572 385960 14600
rect 154632 14560 154638 14572
rect 385954 14560 385960 14572
rect 386012 14560 386018 14612
rect 114002 14492 114008 14544
rect 114060 14532 114066 14544
rect 134150 14532 134156 14544
rect 114060 14504 134156 14532
rect 114060 14492 114066 14504
rect 134150 14492 134156 14504
rect 134208 14492 134214 14544
rect 158898 14492 158904 14544
rect 158956 14532 158962 14544
rect 436738 14532 436744 14544
rect 158956 14504 436744 14532
rect 158956 14492 158962 14504
rect 436738 14492 436744 14504
rect 436796 14492 436802 14544
rect 39114 14424 39120 14476
rect 39172 14464 39178 14476
rect 120718 14464 120724 14476
rect 39172 14436 120724 14464
rect 39172 14424 39178 14436
rect 120718 14424 120724 14436
rect 120776 14424 120782 14476
rect 164326 14424 164332 14476
rect 164384 14464 164390 14476
rect 502978 14464 502984 14476
rect 164384 14436 502984 14464
rect 164384 14424 164390 14436
rect 502978 14424 502984 14436
rect 503036 14424 503042 14476
rect 151998 13404 152004 13456
rect 152056 13444 152062 13456
rect 345290 13444 345296 13456
rect 152056 13416 345296 13444
rect 152056 13404 152062 13416
rect 345290 13404 345296 13416
rect 345348 13404 345354 13456
rect 151906 13336 151912 13388
rect 151964 13376 151970 13388
rect 349154 13376 349160 13388
rect 151964 13348 349160 13376
rect 151964 13336 151970 13348
rect 349154 13336 349160 13348
rect 349212 13336 349218 13388
rect 153378 13268 153384 13320
rect 153436 13308 153442 13320
rect 365714 13308 365720 13320
rect 153436 13280 365720 13308
rect 153436 13268 153442 13280
rect 365714 13268 365720 13280
rect 365772 13268 365778 13320
rect 157610 13200 157616 13252
rect 157668 13240 157674 13252
rect 417418 13240 417424 13252
rect 157668 13212 417424 13240
rect 157668 13200 157674 13212
rect 417418 13200 417424 13212
rect 417476 13200 417482 13252
rect 158806 13132 158812 13184
rect 158864 13172 158870 13184
rect 429194 13172 429200 13184
rect 158864 13144 429200 13172
rect 158864 13132 158870 13144
rect 429194 13132 429200 13144
rect 429252 13132 429258 13184
rect 160186 13064 160192 13116
rect 160244 13104 160250 13116
rect 453298 13104 453304 13116
rect 160244 13076 453304 13104
rect 160244 13064 160250 13076
rect 453298 13064 453304 13076
rect 453356 13064 453362 13116
rect 143626 11976 143632 12028
rect 143684 12016 143690 12028
rect 237650 12016 237656 12028
rect 143684 11988 237656 12016
rect 143684 11976 143690 11988
rect 237650 11976 237656 11988
rect 237708 11976 237714 12028
rect 150342 11908 150348 11960
rect 150400 11948 150406 11960
rect 313826 11948 313832 11960
rect 150400 11920 313832 11948
rect 150400 11908 150406 11920
rect 313826 11908 313832 11920
rect 313884 11908 313890 11960
rect 135806 11840 135812 11892
rect 135864 11840 135870 11892
rect 157426 11840 157432 11892
rect 157484 11880 157490 11892
rect 414290 11880 414296 11892
rect 157484 11852 414296 11880
rect 157484 11840 157490 11852
rect 414290 11840 414296 11852
rect 414348 11840 414354 11892
rect 135714 11636 135720 11688
rect 135772 11676 135778 11688
rect 135824 11676 135852 11840
rect 157518 11772 157524 11824
rect 157576 11812 157582 11824
rect 415486 11812 415492 11824
rect 157576 11784 415492 11812
rect 157576 11772 157582 11784
rect 415486 11772 415492 11784
rect 415544 11772 415550 11824
rect 165798 11704 165804 11756
rect 165856 11744 165862 11756
rect 523770 11744 523776 11756
rect 165856 11716 523776 11744
rect 165856 11704 165862 11716
rect 523770 11704 523776 11716
rect 523828 11704 523834 11756
rect 135772 11648 135852 11676
rect 135772 11636 135778 11648
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 184934 11636 184940 11688
rect 184992 11676 184998 11688
rect 186130 11676 186136 11688
rect 184992 11648 186136 11676
rect 184992 11636 184998 11648
rect 186130 11636 186136 11648
rect 186188 11636 186194 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 106458 10616 106464 10668
rect 106516 10656 106522 10668
rect 132954 10656 132960 10668
rect 106516 10628 132960 10656
rect 106516 10616 106522 10628
rect 132954 10616 132960 10628
rect 133012 10616 133018 10668
rect 99834 10548 99840 10600
rect 99892 10588 99898 10600
rect 133046 10588 133052 10600
rect 99892 10560 133052 10588
rect 99892 10548 99898 10560
rect 133046 10548 133052 10560
rect 133104 10548 133110 10600
rect 147674 10548 147680 10600
rect 147732 10588 147738 10600
rect 295610 10588 295616 10600
rect 147732 10560 295616 10588
rect 147732 10548 147738 10560
rect 295610 10548 295616 10560
rect 295668 10548 295674 10600
rect 81618 10480 81624 10532
rect 81676 10520 81682 10532
rect 131574 10520 131580 10532
rect 81676 10492 131580 10520
rect 81676 10480 81682 10492
rect 131574 10480 131580 10492
rect 131632 10480 131638 10532
rect 154482 10480 154488 10532
rect 154540 10520 154546 10532
rect 364610 10520 364616 10532
rect 154540 10492 364616 10520
rect 154540 10480 154546 10492
rect 364610 10480 364616 10492
rect 364668 10480 364674 10532
rect 35986 10412 35992 10464
rect 36044 10452 36050 10464
rect 127250 10452 127256 10464
rect 36044 10424 127256 10452
rect 36044 10412 36050 10424
rect 127250 10412 127256 10424
rect 127308 10412 127314 10464
rect 156046 10412 156052 10464
rect 156104 10452 156110 10464
rect 394234 10452 394240 10464
rect 156104 10424 394240 10452
rect 156104 10412 156110 10424
rect 394234 10412 394240 10424
rect 394292 10412 394298 10464
rect 28442 10344 28448 10396
rect 28500 10384 28506 10396
rect 127158 10384 127164 10396
rect 28500 10356 127164 10384
rect 28500 10344 28506 10356
rect 127158 10344 127164 10356
rect 127216 10344 127222 10396
rect 156138 10344 156144 10396
rect 156196 10384 156202 10396
rect 398926 10384 398932 10396
rect 156196 10356 398932 10384
rect 156196 10344 156202 10356
rect 398926 10344 398932 10356
rect 398984 10344 398990 10396
rect 11146 10276 11152 10328
rect 11204 10316 11210 10328
rect 126146 10316 126152 10328
rect 11204 10288 126152 10316
rect 11204 10276 11210 10288
rect 126146 10276 126152 10288
rect 126204 10276 126210 10328
rect 163130 10276 163136 10328
rect 163188 10316 163194 10328
rect 486418 10316 486424 10328
rect 163188 10288 486424 10316
rect 163188 10276 163194 10288
rect 486418 10276 486424 10288
rect 486476 10276 486482 10328
rect 67910 9324 67916 9376
rect 67968 9364 67974 9376
rect 130194 9364 130200 9376
rect 67968 9336 130200 9364
rect 67968 9324 67974 9336
rect 130194 9324 130200 9336
rect 130252 9324 130258 9376
rect 64322 9256 64328 9308
rect 64380 9296 64386 9308
rect 126330 9296 126336 9308
rect 64380 9268 126336 9296
rect 64380 9256 64386 9268
rect 126330 9256 126336 9268
rect 126388 9256 126394 9308
rect 144914 9256 144920 9308
rect 144972 9296 144978 9308
rect 260650 9296 260656 9308
rect 144972 9268 260656 9296
rect 144972 9256 144978 9268
rect 260650 9256 260656 9268
rect 260708 9256 260714 9308
rect 63218 9188 63224 9240
rect 63276 9228 63282 9240
rect 130102 9228 130108 9240
rect 63276 9200 130108 9228
rect 63276 9188 63282 9200
rect 130102 9188 130108 9200
rect 130160 9188 130166 9240
rect 146294 9188 146300 9240
rect 146352 9228 146358 9240
rect 278314 9228 278320 9240
rect 146352 9200 278320 9228
rect 146352 9188 146358 9200
rect 278314 9188 278320 9200
rect 278372 9188 278378 9240
rect 60826 9120 60832 9172
rect 60884 9160 60890 9172
rect 129090 9160 129096 9172
rect 60884 9132 129096 9160
rect 60884 9120 60890 9132
rect 129090 9120 129096 9132
rect 129148 9120 129154 9172
rect 151814 9120 151820 9172
rect 151872 9160 151878 9172
rect 343358 9160 343364 9172
rect 151872 9132 343364 9160
rect 151872 9120 151878 9132
rect 343358 9120 343364 9132
rect 343416 9120 343422 9172
rect 53742 9052 53748 9104
rect 53800 9092 53806 9104
rect 128722 9092 128728 9104
rect 53800 9064 128728 9092
rect 53800 9052 53806 9064
rect 128722 9052 128728 9064
rect 128780 9052 128786 9104
rect 161658 9052 161664 9104
rect 161716 9092 161722 9104
rect 471054 9092 471060 9104
rect 161716 9064 471060 9092
rect 161716 9052 161722 9064
rect 471054 9052 471060 9064
rect 471112 9052 471118 9104
rect 50154 8984 50160 9036
rect 50212 9024 50218 9036
rect 126974 9024 126980 9036
rect 50212 8996 126980 9024
rect 50212 8984 50218 8996
rect 126974 8984 126980 8996
rect 127032 8984 127038 9036
rect 163038 8984 163044 9036
rect 163096 9024 163102 9036
rect 492306 9024 492312 9036
rect 163096 8996 492312 9024
rect 163096 8984 163102 8996
rect 492306 8984 492312 8996
rect 492364 8984 492370 9036
rect 566 8916 572 8968
rect 624 8956 630 8968
rect 124214 8956 124220 8968
rect 624 8928 124220 8956
rect 624 8916 630 8928
rect 124214 8916 124220 8928
rect 124272 8916 124278 8968
rect 169938 8916 169944 8968
rect 169996 8956 170002 8968
rect 571518 8956 571524 8968
rect 169996 8928 571524 8956
rect 169996 8916 170002 8928
rect 571518 8916 571524 8928
rect 571576 8916 571582 8968
rect 116394 7896 116400 7948
rect 116452 7936 116458 7948
rect 134058 7936 134064 7948
rect 116452 7908 134064 7936
rect 116452 7896 116458 7908
rect 134058 7896 134064 7908
rect 134116 7896 134122 7948
rect 142246 7896 142252 7948
rect 142304 7936 142310 7948
rect 225138 7936 225144 7948
rect 142304 7908 225144 7936
rect 142304 7896 142310 7908
rect 225138 7896 225144 7908
rect 225196 7896 225202 7948
rect 105722 7828 105728 7880
rect 105780 7868 105786 7880
rect 132862 7868 132868 7880
rect 105780 7840 132868 7868
rect 105780 7828 105786 7840
rect 132862 7828 132868 7840
rect 132920 7828 132926 7880
rect 143534 7828 143540 7880
rect 143592 7868 143598 7880
rect 242986 7868 242992 7880
rect 143592 7840 242992 7868
rect 143592 7828 143598 7840
rect 242986 7828 242992 7840
rect 243044 7828 243050 7880
rect 98638 7760 98644 7812
rect 98696 7800 98702 7812
rect 132770 7800 132776 7812
rect 98696 7772 132776 7800
rect 98696 7760 98702 7772
rect 132770 7760 132776 7772
rect 132828 7760 132834 7812
rect 155954 7760 155960 7812
rect 156012 7800 156018 7812
rect 401318 7800 401324 7812
rect 156012 7772 401324 7800
rect 156012 7760 156018 7772
rect 401318 7760 401324 7772
rect 401376 7760 401382 7812
rect 48958 7692 48964 7744
rect 49016 7732 49022 7744
rect 128630 7732 128636 7744
rect 49016 7704 128636 7732
rect 49016 7692 49022 7704
rect 128630 7692 128636 7704
rect 128688 7692 128694 7744
rect 160094 7692 160100 7744
rect 160152 7732 160158 7744
rect 446214 7732 446220 7744
rect 160152 7704 446220 7732
rect 160152 7692 160158 7704
rect 446214 7692 446220 7704
rect 446272 7692 446278 7744
rect 44266 7624 44272 7676
rect 44324 7664 44330 7676
rect 128538 7664 128544 7676
rect 44324 7636 128544 7664
rect 44324 7624 44330 7636
rect 128538 7624 128544 7636
rect 128596 7624 128602 7676
rect 161566 7624 161572 7676
rect 161624 7664 161630 7676
rect 469858 7664 469864 7676
rect 161624 7636 469864 7664
rect 161624 7624 161630 7636
rect 469858 7624 469864 7636
rect 469916 7624 469922 7676
rect 9950 7556 9956 7608
rect 10008 7596 10014 7608
rect 126054 7596 126060 7608
rect 10008 7568 126060 7596
rect 10008 7556 10014 7568
rect 126054 7556 126060 7568
rect 126112 7556 126118 7608
rect 164234 7556 164240 7608
rect 164292 7596 164298 7608
rect 504174 7596 504180 7608
rect 164292 7568 504180 7596
rect 164292 7556 164298 7568
rect 504174 7556 504180 7568
rect 504232 7556 504238 7608
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 151078 6740 151084 6792
rect 151136 6780 151142 6792
rect 323302 6780 323308 6792
rect 151136 6752 323308 6780
rect 151136 6740 151142 6752
rect 323302 6740 323308 6752
rect 323360 6740 323366 6792
rect 150894 6672 150900 6724
rect 150952 6712 150958 6724
rect 326798 6712 326804 6724
rect 150952 6684 326804 6712
rect 150952 6672 150958 6684
rect 326798 6672 326804 6684
rect 326856 6672 326862 6724
rect 115198 6604 115204 6656
rect 115256 6644 115262 6656
rect 134702 6644 134708 6656
rect 115256 6616 134708 6644
rect 115256 6604 115262 6616
rect 134702 6604 134708 6616
rect 134760 6604 134766 6656
rect 150986 6604 150992 6656
rect 151044 6644 151050 6656
rect 329190 6644 329196 6656
rect 151044 6616 329196 6644
rect 151044 6604 151050 6616
rect 329190 6604 329196 6616
rect 329248 6604 329254 6656
rect 104526 6536 104532 6588
rect 104584 6576 104590 6588
rect 132678 6576 132684 6588
rect 104584 6548 132684 6576
rect 104584 6536 104590 6548
rect 132678 6536 132684 6548
rect 132736 6536 132742 6588
rect 150802 6536 150808 6588
rect 150860 6576 150866 6588
rect 330386 6576 330392 6588
rect 150860 6548 330392 6576
rect 150860 6536 150866 6548
rect 330386 6536 330392 6548
rect 330444 6536 330450 6588
rect 84470 6468 84476 6520
rect 84528 6508 84534 6520
rect 131298 6508 131304 6520
rect 84528 6480 131304 6508
rect 84528 6468 84534 6480
rect 131298 6468 131304 6480
rect 131356 6468 131362 6520
rect 157334 6468 157340 6520
rect 157392 6508 157398 6520
rect 410794 6508 410800 6520
rect 157392 6480 410800 6508
rect 157392 6468 157398 6480
rect 410794 6468 410800 6480
rect 410852 6468 410858 6520
rect 80882 6400 80888 6452
rect 80940 6440 80946 6452
rect 131482 6440 131488 6452
rect 80940 6412 131488 6440
rect 80940 6400 80946 6412
rect 131482 6400 131488 6412
rect 131540 6400 131546 6452
rect 175918 6400 175924 6452
rect 175976 6440 175982 6452
rect 433242 6440 433248 6452
rect 175976 6412 433248 6440
rect 175976 6400 175982 6412
rect 433242 6400 433248 6412
rect 433300 6400 433306 6452
rect 77386 6332 77392 6384
rect 77444 6372 77450 6384
rect 131390 6372 131396 6384
rect 77444 6344 131396 6372
rect 77444 6332 77450 6344
rect 131390 6332 131396 6344
rect 131448 6332 131454 6384
rect 158714 6332 158720 6384
rect 158772 6372 158778 6384
rect 441522 6372 441528 6384
rect 158772 6344 441528 6372
rect 158772 6332 158778 6344
rect 441522 6332 441528 6344
rect 441580 6332 441586 6384
rect 25314 6264 25320 6316
rect 25372 6304 25378 6316
rect 57238 6304 57244 6316
rect 25372 6276 57244 6304
rect 25372 6264 25378 6276
rect 57238 6264 57244 6276
rect 57296 6264 57302 6316
rect 66714 6264 66720 6316
rect 66772 6304 66778 6316
rect 130010 6304 130016 6316
rect 66772 6276 130016 6304
rect 66772 6264 66778 6276
rect 130010 6264 130016 6276
rect 130068 6264 130074 6316
rect 161474 6264 161480 6316
rect 161532 6304 161538 6316
rect 467466 6304 467472 6316
rect 161532 6276 467472 6304
rect 161532 6264 161538 6276
rect 467466 6264 467472 6276
rect 467524 6264 467530 6316
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 127526 6236 127532 6248
rect 33652 6208 127532 6236
rect 33652 6196 33658 6208
rect 127526 6196 127532 6208
rect 127584 6196 127590 6248
rect 140406 6196 140412 6248
rect 140464 6236 140470 6248
rect 156598 6236 156604 6248
rect 140464 6208 156604 6236
rect 140464 6196 140470 6208
rect 156598 6196 156604 6208
rect 156656 6196 156662 6248
rect 169846 6196 169852 6248
rect 169904 6236 169910 6248
rect 572714 6236 572720 6248
rect 169904 6208 572720 6236
rect 169904 6196 169910 6208
rect 572714 6196 572720 6208
rect 572772 6196 572778 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 125962 6168 125968 6180
rect 18288 6140 125968 6168
rect 18288 6128 18294 6140
rect 125962 6128 125968 6140
rect 126020 6128 126026 6180
rect 138290 6128 138296 6180
rect 138348 6168 138354 6180
rect 162486 6168 162492 6180
rect 138348 6140 162492 6168
rect 138348 6128 138354 6140
rect 162486 6128 162492 6140
rect 162544 6128 162550 6180
rect 169754 6128 169760 6180
rect 169812 6168 169818 6180
rect 576302 6168 576308 6180
rect 169812 6140 576308 6168
rect 169812 6128 169818 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 101030 5312 101036 5364
rect 101088 5352 101094 5364
rect 133138 5352 133144 5364
rect 101088 5324 133144 5352
rect 101088 5312 101094 5324
rect 133138 5312 133144 5324
rect 133196 5312 133202 5364
rect 97442 5244 97448 5296
rect 97500 5284 97506 5296
rect 132586 5284 132592 5296
rect 97500 5256 132592 5284
rect 97500 5244 97506 5256
rect 132586 5244 132592 5256
rect 132644 5244 132650 5296
rect 86862 5176 86868 5228
rect 86920 5216 86926 5228
rect 132034 5216 132040 5228
rect 86920 5188 132040 5216
rect 86920 5176 86926 5188
rect 132034 5176 132040 5188
rect 132092 5176 132098 5228
rect 138106 5176 138112 5228
rect 138164 5216 138170 5228
rect 169570 5216 169576 5228
rect 138164 5188 169576 5216
rect 138164 5176 138170 5188
rect 169570 5176 169576 5188
rect 169628 5176 169634 5228
rect 28966 5120 38654 5148
rect 15930 5040 15936 5092
rect 15988 5080 15994 5092
rect 28966 5080 28994 5120
rect 15988 5052 28994 5080
rect 38626 5080 38654 5120
rect 59630 5108 59636 5160
rect 59688 5148 59694 5160
rect 129918 5148 129924 5160
rect 59688 5120 129924 5148
rect 59688 5108 59694 5120
rect 129918 5108 129924 5120
rect 129976 5108 129982 5160
rect 142154 5108 142160 5160
rect 142212 5148 142218 5160
rect 220446 5148 220452 5160
rect 142212 5120 220452 5148
rect 142212 5108 142218 5120
rect 220446 5108 220452 5120
rect 220504 5108 220510 5160
rect 46198 5080 46204 5092
rect 38626 5052 46204 5080
rect 15988 5040 15994 5052
rect 46198 5040 46204 5052
rect 46256 5040 46262 5092
rect 52546 5040 52552 5092
rect 52604 5080 52610 5092
rect 129642 5080 129648 5092
rect 52604 5052 129648 5080
rect 52604 5040 52610 5052
rect 129642 5040 129648 5052
rect 129700 5040 129706 5092
rect 137094 5040 137100 5092
rect 137152 5080 137158 5092
rect 148318 5080 148324 5092
rect 137152 5052 148324 5080
rect 137152 5040 137158 5052
rect 148318 5040 148324 5052
rect 148376 5040 148382 5092
rect 153286 5040 153292 5092
rect 153344 5080 153350 5092
rect 365806 5080 365812 5092
rect 153344 5052 365812 5080
rect 153344 5040 153350 5052
rect 365806 5040 365812 5052
rect 365864 5040 365870 5092
rect 33226 4972 33232 5024
rect 33284 5012 33290 5024
rect 127434 5012 127440 5024
rect 33284 4984 127440 5012
rect 33284 4972 33290 4984
rect 127434 4972 127440 4984
rect 127492 4972 127498 5024
rect 138014 4972 138020 5024
rect 138072 5012 138078 5024
rect 171962 5012 171968 5024
rect 138072 4984 171968 5012
rect 138072 4972 138078 4984
rect 171962 4972 171968 4984
rect 172020 4972 172026 5024
rect 180058 4972 180064 5024
rect 180116 5012 180122 5024
rect 450906 5012 450912 5024
rect 180116 4984 450912 5012
rect 180116 4972 180122 4984
rect 450906 4972 450912 4984
rect 450964 4972 450970 5024
rect 6454 4904 6460 4956
rect 6512 4944 6518 4956
rect 22738 4944 22744 4956
rect 6512 4916 22744 4944
rect 6512 4904 6518 4916
rect 22738 4904 22744 4916
rect 22796 4904 22802 4956
rect 24210 4904 24216 4956
rect 24268 4944 24274 4956
rect 122098 4944 122104 4956
rect 24268 4916 122104 4944
rect 24268 4904 24274 4916
rect 122098 4904 122104 4916
rect 122156 4904 122162 4956
rect 136910 4904 136916 4956
rect 136968 4944 136974 4956
rect 150618 4944 150624 4956
rect 136968 4916 150624 4944
rect 136968 4904 136974 4916
rect 150618 4904 150624 4916
rect 150676 4904 150682 4956
rect 162946 4904 162952 4956
rect 163004 4944 163010 4956
rect 487614 4944 487620 4956
rect 163004 4916 487620 4944
rect 163004 4904 163010 4916
rect 487614 4904 487620 4916
rect 487672 4904 487678 4956
rect 13538 4836 13544 4888
rect 13596 4876 13602 4888
rect 125870 4876 125876 4888
rect 13596 4848 125876 4876
rect 13596 4836 13602 4848
rect 125870 4836 125876 4848
rect 125928 4836 125934 4888
rect 137002 4836 137008 4888
rect 137060 4876 137066 4888
rect 157794 4876 157800 4888
rect 137060 4848 157800 4876
rect 137060 4836 137066 4848
rect 157794 4836 157800 4848
rect 157852 4836 157858 4888
rect 165614 4836 165620 4888
rect 165672 4876 165678 4888
rect 523034 4876 523040 4888
rect 165672 4848 523040 4876
rect 165672 4836 165678 4848
rect 523034 4836 523040 4848
rect 523092 4836 523098 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 125778 4808 125784 4820
rect 8812 4780 125784 4808
rect 8812 4768 8818 4780
rect 125778 4768 125784 4780
rect 125836 4768 125842 4820
rect 138198 4768 138204 4820
rect 138256 4808 138262 4820
rect 164878 4808 164884 4820
rect 138256 4780 164884 4808
rect 138256 4768 138262 4780
rect 164878 4768 164884 4780
rect 164936 4768 164942 4820
rect 165706 4768 165712 4820
rect 165764 4808 165770 4820
rect 527818 4808 527824 4820
rect 165764 4780 527824 4808
rect 165764 4768 165770 4780
rect 527818 4768 527824 4780
rect 527876 4768 527882 4820
rect 138934 4360 138940 4412
rect 138992 4400 138998 4412
rect 143534 4400 143540 4412
rect 138992 4372 143540 4400
rect 138992 4360 138998 4372
rect 143534 4360 143540 4372
rect 143592 4360 143598 4412
rect 242894 4156 242900 4208
rect 242952 4196 242958 4208
rect 244090 4196 244096 4208
rect 242952 4168 244096 4196
rect 242952 4156 242958 4168
rect 244090 4156 244096 4168
rect 244148 4156 244154 4208
rect 251174 4156 251180 4208
rect 251232 4196 251238 4208
rect 252370 4196 252376 4208
rect 251232 4168 252376 4196
rect 251232 4156 251238 4168
rect 252370 4156 252376 4168
rect 252428 4156 252434 4208
rect 276014 4156 276020 4208
rect 276072 4196 276078 4208
rect 276750 4196 276756 4208
rect 276072 4168 276756 4196
rect 276072 4156 276078 4168
rect 276750 4156 276756 4168
rect 276808 4156 276814 4208
rect 119890 4088 119896 4140
rect 119948 4128 119954 4140
rect 124858 4128 124864 4140
rect 119948 4100 124864 4128
rect 119948 4088 119954 4100
rect 124858 4088 124864 4100
rect 124916 4088 124922 4140
rect 125870 4088 125876 4140
rect 125928 4128 125934 4140
rect 134518 4128 134524 4140
rect 125928 4100 134524 4128
rect 125928 4088 125934 4100
rect 134518 4088 134524 4100
rect 134576 4088 134582 4140
rect 151538 4088 151544 4140
rect 151596 4128 151602 4140
rect 325602 4128 325608 4140
rect 151596 4100 325608 4128
rect 151596 4088 151602 4100
rect 325602 4088 325608 4100
rect 325660 4088 325666 4140
rect 138658 4020 138664 4072
rect 138716 4060 138722 4072
rect 145926 4060 145932 4072
rect 138716 4032 145932 4060
rect 138716 4020 138722 4032
rect 145926 4020 145932 4032
rect 145984 4020 145990 4072
rect 150526 4020 150532 4072
rect 150584 4060 150590 4072
rect 327994 4060 328000 4072
rect 150584 4032 328000 4060
rect 150584 4020 150590 4032
rect 327994 4020 328000 4032
rect 328052 4020 328058 4072
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 126606 3992 126612 4004
rect 12400 3964 126612 3992
rect 12400 3952 12406 3964
rect 126606 3952 126612 3964
rect 126664 3952 126670 4004
rect 135806 3952 135812 4004
rect 135864 3992 135870 4004
rect 141234 3992 141240 4004
rect 135864 3964 141240 3992
rect 135864 3952 135870 3964
rect 141234 3952 141240 3964
rect 141292 3952 141298 4004
rect 150894 3952 150900 4004
rect 150952 3992 150958 4004
rect 331582 3992 331588 4004
rect 150952 3964 331588 3992
rect 150952 3952 150958 3964
rect 331582 3952 331588 3964
rect 331640 3952 331646 4004
rect 137738 3884 137744 3936
rect 137796 3924 137802 3936
rect 144730 3924 144736 3936
rect 137796 3896 144736 3924
rect 137796 3884 137802 3896
rect 144730 3884 144736 3896
rect 144788 3884 144794 3936
rect 172146 3884 172152 3936
rect 172204 3924 172210 3936
rect 356330 3924 356336 3936
rect 172204 3896 356336 3924
rect 172204 3884 172210 3896
rect 356330 3884 356336 3896
rect 356388 3884 356394 3936
rect 467098 3884 467104 3936
rect 467156 3924 467162 3936
rect 534902 3924 534908 3936
rect 467156 3896 534908 3924
rect 467156 3884 467162 3896
rect 534902 3884 534908 3896
rect 534960 3884 534966 3936
rect 83274 3816 83280 3868
rect 83332 3856 83338 3868
rect 131850 3856 131856 3868
rect 83332 3828 131856 3856
rect 83332 3816 83338 3828
rect 131850 3816 131856 3828
rect 131908 3816 131914 3868
rect 135530 3816 135536 3868
rect 135588 3856 135594 3868
rect 138842 3856 138848 3868
rect 135588 3828 138848 3856
rect 135588 3816 135594 3828
rect 138842 3816 138848 3828
rect 138900 3816 138906 3868
rect 142982 3816 142988 3868
rect 143040 3856 143046 3868
rect 151814 3856 151820 3868
rect 143040 3828 151820 3856
rect 143040 3816 143046 3828
rect 151814 3816 151820 3828
rect 151872 3816 151878 3868
rect 172054 3816 172060 3868
rect 172112 3856 172118 3868
rect 303154 3856 303160 3868
rect 172112 3828 303160 3856
rect 172112 3816 172118 3828
rect 303154 3816 303160 3828
rect 303212 3816 303218 3868
rect 319438 3816 319444 3868
rect 319496 3856 319502 3868
rect 583386 3856 583392 3868
rect 319496 3828 583392 3856
rect 319496 3816 319502 3828
rect 583386 3816 583392 3828
rect 583444 3816 583450 3868
rect 76190 3748 76196 3800
rect 76248 3788 76254 3800
rect 128998 3788 129004 3800
rect 76248 3760 129004 3788
rect 76248 3748 76254 3760
rect 128998 3748 129004 3760
rect 129056 3748 129062 3800
rect 131758 3748 131764 3800
rect 131816 3788 131822 3800
rect 135714 3788 135720 3800
rect 131816 3760 135720 3788
rect 131816 3748 131822 3760
rect 135714 3748 135720 3760
rect 135772 3748 135778 3800
rect 136818 3748 136824 3800
rect 136876 3788 136882 3800
rect 136876 3760 137784 3788
rect 136876 3748 136882 3760
rect 69106 3680 69112 3732
rect 69164 3720 69170 3732
rect 130654 3720 130660 3732
rect 69164 3692 130660 3720
rect 69164 3680 69170 3692
rect 130654 3680 130660 3692
rect 130712 3680 130718 3732
rect 135438 3680 135444 3732
rect 135496 3720 135502 3732
rect 137646 3720 137652 3732
rect 135496 3692 137652 3720
rect 135496 3680 135502 3692
rect 137646 3680 137652 3692
rect 137704 3680 137710 3732
rect 137756 3720 137784 3760
rect 140130 3748 140136 3800
rect 140188 3788 140194 3800
rect 149514 3788 149520 3800
rect 140188 3760 149520 3788
rect 140188 3748 140194 3760
rect 149514 3748 149520 3760
rect 149572 3748 149578 3800
rect 152550 3748 152556 3800
rect 152608 3788 152614 3800
rect 168374 3788 168380 3800
rect 152608 3760 168380 3788
rect 152608 3748 152614 3760
rect 168374 3748 168380 3760
rect 168432 3748 168438 3800
rect 178678 3748 178684 3800
rect 178736 3788 178742 3800
rect 475746 3788 475752 3800
rect 178736 3760 475752 3788
rect 178736 3748 178742 3760
rect 475746 3748 475752 3760
rect 475804 3748 475810 3800
rect 154206 3720 154212 3732
rect 137756 3692 154212 3720
rect 154206 3680 154212 3692
rect 154264 3680 154270 3732
rect 163958 3680 163964 3732
rect 164016 3720 164022 3732
rect 491110 3720 491116 3732
rect 164016 3692 491116 3720
rect 164016 3680 164022 3692
rect 491110 3680 491116 3692
rect 491168 3680 491174 3732
rect 62022 3612 62028 3664
rect 62080 3652 62086 3664
rect 122190 3652 122196 3664
rect 62080 3624 122196 3652
rect 62080 3612 62086 3624
rect 122190 3612 122196 3624
rect 122248 3612 122254 3664
rect 127618 3652 127624 3664
rect 122806 3624 127624 3652
rect 47854 3544 47860 3596
rect 47912 3584 47918 3596
rect 122806 3584 122834 3624
rect 127618 3612 127624 3624
rect 127676 3612 127682 3664
rect 132954 3612 132960 3664
rect 133012 3652 133018 3664
rect 135622 3652 135628 3664
rect 133012 3624 135628 3652
rect 133012 3612 133018 3624
rect 135622 3612 135628 3624
rect 135680 3612 135686 3664
rect 135898 3612 135904 3664
rect 135956 3652 135962 3664
rect 140038 3652 140044 3664
rect 135956 3624 140044 3652
rect 135956 3612 135962 3624
rect 140038 3612 140044 3624
rect 140096 3612 140102 3664
rect 155402 3652 155408 3664
rect 140148 3624 155408 3652
rect 47912 3556 122834 3584
rect 47912 3544 47918 3556
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 130378 3584 130384 3596
rect 127032 3556 130384 3584
rect 127032 3544 127038 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 135346 3544 135352 3596
rect 135404 3584 135410 3596
rect 136450 3584 136456 3596
rect 135404 3556 136456 3584
rect 135404 3544 135410 3556
rect 136450 3544 136456 3556
rect 136508 3544 136514 3596
rect 136726 3544 136732 3596
rect 136784 3584 136790 3596
rect 140148 3584 140176 3624
rect 155402 3612 155408 3624
rect 155460 3612 155466 3664
rect 171870 3612 171876 3664
rect 171928 3652 171934 3664
rect 501782 3652 501788 3664
rect 171928 3624 501788 3652
rect 171928 3612 171934 3624
rect 501782 3612 501788 3624
rect 501840 3612 501846 3664
rect 147122 3584 147128 3596
rect 136784 3556 140176 3584
rect 140240 3556 147128 3584
rect 136784 3544 136790 3556
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 126422 3516 126428 3528
rect 17092 3488 126428 3516
rect 17092 3476 17098 3488
rect 126422 3476 126428 3488
rect 126480 3476 126486 3528
rect 133782 3476 133788 3528
rect 133840 3516 133846 3528
rect 140240 3516 140268 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 147214 3544 147220 3596
rect 147272 3584 147278 3596
rect 167178 3584 167184 3596
rect 147272 3556 167184 3584
rect 147272 3544 147278 3556
rect 167178 3544 167184 3556
rect 167236 3544 167242 3596
rect 171778 3544 171784 3596
rect 171836 3584 171842 3596
rect 515950 3584 515956 3596
rect 171836 3556 515956 3584
rect 171836 3544 171842 3556
rect 515950 3544 515956 3556
rect 516008 3544 516014 3596
rect 133840 3488 140268 3516
rect 133840 3476 133846 3488
rect 141510 3476 141516 3528
rect 141568 3516 141574 3528
rect 166074 3516 166080 3528
rect 141568 3488 166080 3516
rect 141568 3476 141574 3488
rect 166074 3476 166080 3488
rect 166132 3476 166138 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173216 3488 531176 3516
rect 173216 3476 173222 3488
rect 93854 3408 93860 3460
rect 93912 3448 93918 3460
rect 94774 3448 94780 3460
rect 93912 3420 94780 3448
rect 93912 3408 93918 3420
rect 94774 3408 94780 3420
rect 94832 3408 94838 3460
rect 142798 3408 142804 3460
rect 142856 3448 142862 3460
rect 170766 3448 170772 3460
rect 142856 3420 170772 3448
rect 142856 3408 142862 3420
rect 170766 3408 170772 3420
rect 170824 3408 170830 3460
rect 173342 3408 173348 3460
rect 173400 3448 173406 3460
rect 531148 3448 531176 3488
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 533706 3448 533712 3460
rect 173400 3420 528554 3448
rect 531148 3420 533712 3448
rect 173400 3408 173406 3420
rect 150802 3340 150808 3392
rect 150860 3380 150866 3392
rect 322106 3380 322112 3392
rect 150860 3352 322112 3380
rect 150860 3340 150866 3352
rect 322106 3340 322112 3352
rect 322164 3340 322170 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 506474 3340 506480 3392
rect 506532 3380 506538 3392
rect 507302 3380 507308 3392
rect 506532 3352 507308 3380
rect 506532 3340 506538 3352
rect 507302 3340 507308 3352
rect 507360 3340 507366 3392
rect 528526 3380 528554 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 537202 3380 537208 3392
rect 528526 3352 537208 3380
rect 537202 3340 537208 3352
rect 537260 3340 537266 3392
rect 144454 3272 144460 3324
rect 144512 3312 144518 3324
rect 153010 3312 153016 3324
rect 144512 3284 153016 3312
rect 144512 3272 144518 3284
rect 153010 3272 153016 3284
rect 153068 3272 153074 3324
rect 173250 3272 173256 3324
rect 173308 3312 173314 3324
rect 212166 3312 212172 3324
rect 173308 3284 212172 3312
rect 173308 3272 173314 3284
rect 212166 3272 212172 3284
rect 212224 3272 212230 3324
rect 362310 3312 362316 3324
rect 219406 3284 362316 3312
rect 211798 3204 211804 3256
rect 211856 3244 211862 3256
rect 219406 3244 219434 3284
rect 362310 3272 362316 3284
rect 362368 3272 362374 3324
rect 211856 3216 219434 3244
rect 211856 3204 211862 3216
rect 307754 3204 307760 3256
rect 307812 3244 307818 3256
rect 309042 3244 309048 3256
rect 307812 3216 309048 3244
rect 307812 3204 307818 3216
rect 309042 3204 309048 3216
rect 309100 3204 309106 3256
rect 316034 3204 316040 3256
rect 316092 3244 316098 3256
rect 317322 3244 317328 3256
rect 316092 3216 317328 3244
rect 316092 3204 316098 3216
rect 317322 3204 317328 3216
rect 317380 3204 317386 3256
rect 390554 1232 390560 1284
rect 390612 1272 390618 1284
rect 391842 1272 391848 1284
rect 390612 1244 391848 1272
rect 390612 1232 390618 1244
rect 391842 1232 391848 1244
rect 391900 1232 391906 1284
rect 30098 1096 30104 1148
rect 30156 1136 30162 1148
rect 33226 1136 33232 1148
rect 30156 1108 33232 1136
rect 30156 1096 30162 1108
rect 33226 1096 33232 1108
rect 33284 1096 33290 1148
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 410524 700408 410576 700460
rect 429844 700408 429896 700460
rect 409144 700340 409196 700392
rect 494796 700340 494848 700392
rect 364984 700272 365036 700324
rect 374644 700272 374696 700324
rect 407764 700272 407816 700324
rect 559656 700272 559708 700324
rect 332508 699796 332560 699848
rect 334624 699796 334676 699848
rect 150440 699660 150492 699712
rect 154120 699660 154172 699712
rect 195980 699660 196032 699712
rect 202788 699660 202840 699712
rect 231860 699660 231912 699712
rect 235172 699660 235224 699712
rect 348792 699660 348844 699712
rect 350540 699660 350592 699712
rect 281540 698300 281592 698352
rect 283840 698300 283892 698352
rect 300124 698096 300176 698148
rect 302884 698096 302936 698148
rect 350540 698028 350592 698080
rect 353944 698028 353996 698080
rect 229744 695240 229796 695292
rect 231860 695240 231912 695292
rect 280804 694968 280856 695020
rect 281540 694968 281592 695020
rect 189080 694764 189132 694816
rect 195980 694764 196032 694816
rect 258080 694220 258132 694272
rect 267648 694220 267700 694272
rect 149796 693472 149848 693524
rect 150440 693472 150492 693524
rect 302884 692044 302936 692096
rect 313924 692044 313976 692096
rect 374644 691092 374696 691144
rect 377404 691092 377456 691144
rect 247684 689256 247736 689308
rect 258080 689256 258132 689308
rect 181444 688644 181496 688696
rect 189080 688644 189132 688696
rect 206284 687896 206336 687948
rect 218060 687896 218112 687948
rect 148324 687488 148376 687540
rect 149796 687488 149848 687540
rect 334624 686468 334676 686520
rect 349804 686468 349856 686520
rect 221464 685108 221516 685160
rect 229744 685108 229796 685160
rect 353944 683748 353996 683800
rect 358360 683748 358412 683800
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 313924 682388 313976 682440
rect 333244 682388 333296 682440
rect 204260 681708 204312 681760
rect 206284 681708 206336 681760
rect 144184 678920 144236 678972
rect 148324 678988 148376 679040
rect 358360 678444 358412 678496
rect 360844 678444 360896 678496
rect 377404 678240 377456 678292
rect 396448 678240 396500 678292
rect 202144 677016 202196 677068
rect 204260 677016 204312 677068
rect 167000 671304 167052 671356
rect 181444 671304 181496 671356
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 406384 670692 406436 670744
rect 580172 670692 580224 670744
rect 215944 668584 215996 668636
rect 221464 668584 221516 668636
rect 360844 668584 360896 668636
rect 363604 668584 363656 668636
rect 160744 667156 160796 667208
rect 167000 667156 167052 667208
rect 200120 666340 200172 666392
rect 202144 666340 202196 666392
rect 279424 665116 279476 665168
rect 280804 665116 280856 665168
rect 363604 663008 363656 663060
rect 369124 663008 369176 663060
rect 141424 662396 141476 662448
rect 144184 662396 144236 662448
rect 153844 661036 153896 661088
rect 160744 661036 160796 661088
rect 369124 660288 369176 660340
rect 387340 660288 387392 660340
rect 195152 659200 195204 659252
rect 200120 659200 200172 659252
rect 241980 658928 242032 658980
rect 247684 658928 247736 658980
rect 349804 658180 349856 658232
rect 355784 658180 355836 658232
rect 387340 658180 387392 658232
rect 393964 658180 394016 658232
rect 235264 656140 235316 656192
rect 241980 656140 242032 656192
rect 274640 655528 274692 655580
rect 279424 655528 279476 655580
rect 355784 655460 355836 655512
rect 358728 655460 358780 655512
rect 185584 654780 185636 654832
rect 195152 654780 195204 654832
rect 273904 652740 273956 652792
rect 274640 652740 274692 652792
rect 146944 651992 146996 652044
rect 153844 651992 153896 652044
rect 358728 650632 358780 650684
rect 369124 650632 369176 650684
rect 393964 649884 394016 649936
rect 395344 649884 395396 649936
rect 203524 647844 203576 647896
rect 215944 647844 215996 647896
rect 395344 647164 395396 647216
rect 396540 647164 396592 647216
rect 333244 643696 333296 643748
rect 353944 643696 353996 643748
rect 396724 643084 396776 643136
rect 580172 643084 580224 643136
rect 144184 641724 144236 641776
rect 146944 641724 146996 641776
rect 369124 640500 369176 640552
rect 371884 640500 371936 640552
rect 232504 639412 232556 639464
rect 235264 639412 235316 639464
rect 140044 638188 140096 638240
rect 141424 638188 141476 638240
rect 196624 635468 196676 635520
rect 203524 635468 203576 635520
rect 2780 632068 2832 632120
rect 4896 632068 4948 632120
rect 184204 632068 184256 632120
rect 185584 632068 185636 632120
rect 272616 632068 272668 632120
rect 273904 632068 273956 632120
rect 271144 629688 271196 629740
rect 272616 629688 272668 629740
rect 136364 627852 136416 627904
rect 140044 627920 140096 627972
rect 353944 625812 353996 625864
rect 395344 625812 395396 625864
rect 134524 620304 134576 620356
rect 136364 620304 136416 620356
rect 3516 618264 3568 618316
rect 19984 618264 20036 618316
rect 405004 616836 405056 616888
rect 580172 616836 580224 616888
rect 269396 616768 269448 616820
rect 271144 616768 271196 616820
rect 126244 608744 126296 608796
rect 134524 608744 134576 608796
rect 268384 608744 268436 608796
rect 269396 608744 269448 608796
rect 182824 603100 182876 603152
rect 184204 603100 184256 603152
rect 137744 597524 137796 597576
rect 144184 597524 144236 597576
rect 264244 593512 264296 593564
rect 268384 593512 268436 593564
rect 133144 592016 133196 592068
rect 137744 592016 137796 592068
rect 120724 591268 120776 591320
rect 126244 591268 126296 591320
rect 371884 591268 371936 591320
rect 384304 591268 384356 591320
rect 229744 590316 229796 590368
rect 232504 590316 232556 590368
rect 119344 585148 119396 585200
rect 120724 585148 120776 585200
rect 262864 585148 262916 585200
rect 264244 585148 264296 585200
rect 384304 583516 384356 583568
rect 390560 583516 390612 583568
rect 207664 581612 207716 581664
rect 229744 581612 229796 581664
rect 3516 579640 3568 579692
rect 10324 579640 10376 579692
rect 129740 578212 129792 578264
rect 133144 578212 133196 578264
rect 181444 578144 181496 578196
rect 182824 578144 182876 578196
rect 390560 576852 390612 576904
rect 393964 576852 394016 576904
rect 120724 570596 120776 570648
rect 129740 570596 129792 570648
rect 261484 570596 261536 570648
rect 262864 570596 262916 570648
rect 3056 565836 3108 565888
rect 37924 565836 37976 565888
rect 403624 563048 403676 563100
rect 580172 563048 580224 563100
rect 93492 559512 93544 559564
rect 120724 559512 120776 559564
rect 193864 554752 193916 554804
rect 196624 554752 196676 554804
rect 117964 553392 118016 553444
rect 119344 553392 119396 553444
rect 90364 552508 90416 552560
rect 93492 552508 93544 552560
rect 260196 552100 260248 552152
rect 261484 552100 261536 552152
rect 258816 549992 258868 550044
rect 260196 549992 260248 550044
rect 198004 545708 198056 545760
rect 207664 545708 207716 545760
rect 256700 541968 256752 542020
rect 258816 541968 258868 542020
rect 255964 538840 256016 538892
rect 256700 538840 256752 538892
rect 116584 536800 116636 536852
rect 117964 536800 118016 536852
rect 393964 536392 394016 536444
rect 396632 536392 396684 536444
rect 115204 534080 115256 534132
rect 116584 534080 116636 534132
rect 2964 527144 3016 527196
rect 6184 527144 6236 527196
rect 113824 525784 113876 525836
rect 115204 525784 115256 525836
rect 177304 524356 177356 524408
rect 181444 524424 181496 524476
rect 191104 520208 191156 520260
rect 193864 520208 193916 520260
rect 3332 514768 3384 514820
rect 24124 514768 24176 514820
rect 253940 511776 253992 511828
rect 255964 511776 256016 511828
rect 400864 510620 400916 510672
rect 580172 510620 580224 510672
rect 251824 506472 251876 506524
rect 253940 506472 253992 506524
rect 173164 505112 173216 505164
rect 177304 505112 177356 505164
rect 195244 504364 195296 504416
rect 198004 504364 198056 504416
rect 192484 490016 192536 490068
rect 195244 490016 195296 490068
rect 112536 481652 112588 481704
rect 113824 481652 113876 481704
rect 111064 476076 111116 476128
rect 112536 476076 112588 476128
rect 171784 473016 171836 473068
rect 173164 473016 173216 473068
rect 189080 470568 189132 470620
rect 192484 470568 192536 470620
rect 182824 466420 182876 466472
rect 189080 466420 189132 466472
rect 250168 466420 250220 466472
rect 251824 466420 251876 466472
rect 248420 462952 248472 463004
rect 250168 462952 250220 463004
rect 2780 462544 2832 462596
rect 4988 462544 5040 462596
rect 109684 459552 109736 459604
rect 111064 459552 111116 459604
rect 179420 459552 179472 459604
rect 182824 459552 182876 459604
rect 245752 459552 245804 459604
rect 248420 459552 248472 459604
rect 399484 456764 399536 456816
rect 579988 456764 580040 456816
rect 244924 455404 244976 455456
rect 245752 455404 245804 455456
rect 177304 452548 177356 452600
rect 179420 452548 179472 452600
rect 84200 452072 84252 452124
rect 90364 452072 90416 452124
rect 75184 447788 75236 447840
rect 84200 447788 84252 447840
rect 170404 447040 170456 447092
rect 171784 447040 171836 447092
rect 167000 437384 167052 437436
rect 170404 437452 170456 437504
rect 151084 436704 151136 436756
rect 177304 436704 177356 436756
rect 163596 433236 163648 433288
rect 166908 433304 166960 433356
rect 134708 431196 134760 431248
rect 151084 431196 151136 431248
rect 107660 430584 107712 430636
rect 109684 430584 109736 430636
rect 171508 429836 171560 429888
rect 191104 429836 191156 429888
rect 106188 427116 106240 427168
rect 107660 427116 107712 427168
rect 163504 425688 163556 425740
rect 171508 425688 171560 425740
rect 103520 423240 103572 423292
rect 106188 423240 106240 423292
rect 131764 422288 131816 422340
rect 134708 422288 134760 422340
rect 398104 418140 398156 418192
rect 580080 418140 580132 418192
rect 101404 417664 101456 417716
rect 103520 417664 103572 417716
rect 243544 416712 243596 416764
rect 244924 416712 244976 416764
rect 160744 413992 160796 414044
rect 163596 413992 163648 414044
rect 113180 413244 113232 413296
rect 131764 413244 131816 413296
rect 3240 410456 3292 410508
rect 8944 410456 8996 410508
rect 95332 407736 95384 407788
rect 113180 407736 113232 407788
rect 160836 407056 160888 407108
rect 163504 407056 163556 407108
rect 97448 405628 97500 405680
rect 101404 405696 101456 405748
rect 418804 404336 418856 404388
rect 580080 404336 580132 404388
rect 75276 403588 75328 403640
rect 95332 403588 95384 403640
rect 236644 403588 236696 403640
rect 243544 403588 243596 403640
rect 148324 402228 148376 402280
rect 160836 402228 160888 402280
rect 96068 401616 96120 401668
rect 97448 401616 97500 401668
rect 94504 397808 94556 397860
rect 96068 397808 96120 397860
rect 69664 396720 69716 396772
rect 136640 396720 136692 396772
rect 233884 395972 233936 396024
rect 236644 395972 236696 396024
rect 72424 391960 72476 392012
rect 75184 391960 75236 392012
rect 92480 390736 92532 390788
rect 94504 390736 94556 390788
rect 90088 385704 90140 385756
rect 92480 385704 92532 385756
rect 68284 384956 68336 385008
rect 69664 384956 69716 385008
rect 86224 382236 86276 382288
rect 90088 382236 90140 382288
rect 396816 378156 396868 378208
rect 580080 378156 580132 378208
rect 3240 371220 3292 371272
rect 10416 371220 10468 371272
rect 59268 370472 59320 370524
rect 72424 370472 72476 370524
rect 159364 366732 159416 366784
rect 160744 366732 160796 366784
rect 46940 366324 46992 366376
rect 59268 366324 59320 366376
rect 398196 364352 398248 364404
rect 579804 364352 579856 364404
rect 45100 360952 45152 361004
rect 46940 360952 46992 361004
rect 84844 358980 84896 359032
rect 86224 358980 86276 359032
rect 65432 358776 65484 358828
rect 68284 358776 68336 358828
rect 64144 358096 64196 358148
rect 65432 358096 65484 358148
rect 3240 357416 3292 357468
rect 22744 357416 22796 357468
rect 157984 355988 158036 356040
rect 159364 355988 159416 356040
rect 71872 353268 71924 353320
rect 75276 353268 75328 353320
rect 145564 353268 145616 353320
rect 148324 353268 148376 353320
rect 82360 351840 82412 351892
rect 84844 351908 84896 351960
rect 417424 351908 417476 351960
rect 580080 351908 580132 351960
rect 228364 349800 228416 349852
rect 233884 349800 233936 349852
rect 80704 349120 80756 349172
rect 82360 349120 82412 349172
rect 63868 345652 63920 345704
rect 71872 345652 71924 345704
rect 61384 339192 61436 339244
rect 63868 339192 63920 339244
rect 225604 338036 225656 338088
rect 228364 338036 228416 338088
rect 140412 337356 140464 337408
rect 145564 337356 145616 337408
rect 156696 332596 156748 332648
rect 157984 332596 158036 332648
rect 62856 331848 62908 331900
rect 88340 331848 88392 331900
rect 135904 328856 135956 328908
rect 140412 328856 140464 328908
rect 155224 328040 155276 328092
rect 156696 328040 156748 328092
rect 397000 324300 397052 324352
rect 580080 324300 580132 324352
rect 79508 320152 79560 320204
rect 80704 320152 80756 320204
rect 62764 319404 62816 319456
rect 64144 319404 64196 319456
rect 3240 318792 3292 318844
rect 33784 318792 33836 318844
rect 153844 318724 153896 318776
rect 155224 318724 155276 318776
rect 61476 318384 61528 318436
rect 62856 318384 62908 318436
rect 78128 318316 78180 318368
rect 79508 318316 79560 318368
rect 224224 317364 224276 317416
rect 225604 317364 225656 317416
rect 73160 315256 73212 315308
rect 78128 315256 78180 315308
rect 84844 315256 84896 315308
rect 104900 315256 104952 315308
rect 58624 314644 58676 314696
rect 61384 314644 61436 314696
rect 71044 313284 71096 313336
rect 73160 313284 73212 313336
rect 398288 311856 398340 311908
rect 580080 311856 580132 311908
rect 60004 311176 60056 311228
rect 61476 311176 61528 311228
rect 102784 308388 102836 308440
rect 135904 308388 135956 308440
rect 151084 307708 151136 307760
rect 153844 307776 153896 307828
rect 69664 304988 69716 305040
rect 71044 304988 71096 305040
rect 220820 303560 220872 303612
rect 224224 303628 224276 303680
rect 68284 302200 68336 302252
rect 69664 302200 69716 302252
rect 220084 301112 220136 301164
rect 220820 301112 220872 301164
rect 60832 299412 60884 299464
rect 62764 299412 62816 299464
rect 414664 298120 414716 298172
rect 580080 298120 580132 298172
rect 97724 297372 97776 297424
rect 102784 297372 102836 297424
rect 87604 294584 87656 294636
rect 97724 294584 97776 294636
rect 66260 294176 66312 294228
rect 68284 294176 68336 294228
rect 60096 293972 60148 294024
rect 60832 293972 60884 294024
rect 2780 292612 2832 292664
rect 5080 292612 5132 292664
rect 63500 292612 63552 292664
rect 66260 292612 66312 292664
rect 53840 291796 53892 291848
rect 63500 291796 63552 291848
rect 213828 291116 213880 291168
rect 220084 291184 220136 291236
rect 58716 290368 58768 290420
rect 60004 290368 60056 290420
rect 51816 289756 51868 289808
rect 53840 289824 53892 289876
rect 211160 288872 211212 288924
rect 213828 288872 213880 288924
rect 57244 287648 57296 287700
rect 71780 287648 71832 287700
rect 82820 284928 82872 284980
rect 87604 284928 87656 284980
rect 55588 284248 55640 284300
rect 58716 284316 58768 284368
rect 82084 284248 82136 284300
rect 84844 284316 84896 284368
rect 207020 283976 207072 284028
rect 211160 283976 211212 284028
rect 57980 282888 58032 282940
rect 60096 282888 60148 282940
rect 66904 282140 66956 282192
rect 82820 282140 82872 282192
rect 148324 281256 148376 281308
rect 151084 281256 151136 281308
rect 54208 281120 54260 281172
rect 55588 281120 55640 281172
rect 53288 280780 53340 280832
rect 169760 280780 169812 280832
rect 49700 280168 49752 280220
rect 51816 280168 51868 280220
rect 53104 278808 53156 278860
rect 54208 278808 54260 278860
rect 54484 278740 54536 278792
rect 57888 278740 57940 278792
rect 204168 278264 204220 278316
rect 207020 278264 207072 278316
rect 48964 278128 49016 278180
rect 49700 278128 49752 278180
rect 46940 277992 46992 278044
rect 58624 277992 58676 278044
rect 53840 277312 53892 277364
rect 57244 277380 57296 277432
rect 55864 276632 55916 276684
rect 82084 276632 82136 276684
rect 63500 275068 63552 275120
rect 66904 275068 66956 275120
rect 44916 274660 44968 274712
rect 46940 274660 46992 274712
rect 53196 274660 53248 274712
rect 53840 274660 53892 274712
rect 201500 274660 201552 274712
rect 204168 274660 204220 274712
rect 51724 272008 51776 272060
rect 53104 272008 53156 272060
rect 504364 271872 504416 271924
rect 579804 271872 579856 271924
rect 200764 270920 200816 270972
rect 201500 270920 201552 270972
rect 51080 270444 51132 270496
rect 53288 270444 53340 270496
rect 60556 268608 60608 268660
rect 63500 268608 63552 268660
rect 53196 266432 53248 266484
rect 54484 266432 54536 266484
rect 3056 266364 3108 266416
rect 20076 266364 20128 266416
rect 48320 266296 48372 266348
rect 51080 266364 51132 266416
rect 54208 266364 54260 266416
rect 55864 266364 55916 266416
rect 198004 266364 198056 266416
rect 200764 266364 200816 266416
rect 49700 263576 49752 263628
rect 51724 263576 51776 263628
rect 53288 263576 53340 263628
rect 54208 263576 54260 263628
rect 146944 262896 146996 262948
rect 148324 262896 148376 262948
rect 53380 262828 53432 262880
rect 60556 262828 60608 262880
rect 45744 259224 45796 259276
rect 48228 259224 48280 259276
rect 46940 258544 46992 258596
rect 49700 258544 49752 258596
rect 398380 258068 398432 258120
rect 579988 258068 580040 258120
rect 48228 256776 48280 256828
rect 53380 256776 53432 256828
rect 50436 256640 50488 256692
rect 53288 256708 53340 256760
rect 45560 255280 45612 255332
rect 46940 255280 46992 255332
rect 45008 254260 45060 254312
rect 48228 254260 48280 254312
rect 47584 253988 47636 254040
rect 50436 253988 50488 254040
rect 3148 253920 3200 253972
rect 22836 253920 22888 253972
rect 46940 253920 46992 253972
rect 48964 253920 49016 253972
rect 49056 253920 49108 253972
rect 53196 253920 53248 253972
rect 144276 253920 144328 253972
rect 146944 253920 146996 253972
rect 135904 252832 135956 252884
rect 144276 252832 144328 252884
rect 51816 252560 51868 252612
rect 53104 252560 53156 252612
rect 50344 250656 50396 250708
rect 51816 250656 51868 250708
rect 45192 249772 45244 249824
rect 46940 249772 46992 249824
rect 46572 245624 46624 245676
rect 47584 245624 47636 245676
rect 195980 245624 196032 245676
rect 198004 245624 198056 245676
rect 46940 244264 46992 244316
rect 49056 244264 49108 244316
rect 413284 244264 413336 244316
rect 579988 244264 580040 244316
rect 396540 243516 396592 243568
rect 396908 243516 396960 243568
rect 133604 243040 133656 243092
rect 135904 243040 135956 243092
rect 124128 242156 124180 242208
rect 133604 242156 133656 242208
rect 46848 240796 46900 240848
rect 124128 240796 124180 240848
rect 45652 240728 45704 240780
rect 195980 240728 196032 240780
rect 45836 240524 45888 240576
rect 50344 240524 50396 240576
rect 2780 240184 2832 240236
rect 5172 240184 5224 240236
rect 395344 240048 395396 240100
rect 396540 240048 396592 240100
rect 45284 239844 45336 239896
rect 46572 239844 46624 239896
rect 44824 239776 44876 239828
rect 46848 239776 46900 239828
rect 45468 239708 45520 239760
rect 46756 239708 46808 239760
rect 396540 238824 396592 238876
rect 45376 238756 45428 238808
rect 45652 238756 45704 238808
rect 396540 238688 396592 238740
rect 45744 233112 45796 233164
rect 105820 233112 105872 233164
rect 44824 232976 44876 233028
rect 45652 232976 45704 233028
rect 45468 232364 45520 232416
rect 45744 232364 45796 232416
rect 45836 232364 45888 232416
rect 48320 232364 48372 232416
rect 45376 232296 45428 232348
rect 46848 232296 46900 232348
rect 394700 232092 394752 232144
rect 396540 232092 396592 232144
rect 105820 231956 105872 232008
rect 117964 231956 118016 232008
rect 396540 231956 396592 232008
rect 396908 231956 396960 232008
rect 393964 231820 394016 231872
rect 580080 231820 580132 231872
rect 45744 231752 45796 231804
rect 50620 231752 50672 231804
rect 3332 231140 3384 231192
rect 179420 231140 179472 231192
rect 4068 231072 4120 231124
rect 180800 231072 180852 231124
rect 45284 231004 45336 231056
rect 159364 231004 159416 231056
rect 48320 230936 48372 230988
rect 72424 230936 72476 230988
rect 45192 230460 45244 230512
rect 46940 230460 46992 230512
rect 46848 230392 46900 230444
rect 49608 230392 49660 230444
rect 45652 230324 45704 230376
rect 51540 230324 51592 230376
rect 392676 229780 392728 229832
rect 396632 229780 396684 229832
rect 117964 229712 118016 229764
rect 131764 229712 131816 229764
rect 390928 229508 390980 229560
rect 394700 229508 394752 229560
rect 157984 228420 158036 228472
rect 266544 228420 266596 228472
rect 267004 228420 267056 228472
rect 356520 228420 356572 228472
rect 118792 228352 118844 228404
rect 580724 228352 580776 228404
rect 50620 227808 50672 227860
rect 56508 227808 56560 227860
rect 2872 227740 2924 227792
rect 138664 227740 138716 227792
rect 49700 227468 49752 227520
rect 52368 227468 52420 227520
rect 72424 226992 72476 227044
rect 77944 226992 77996 227044
rect 377312 226992 377364 227044
rect 396540 226992 396592 227044
rect 384396 226856 384448 226908
rect 390928 226856 390980 226908
rect 46940 225564 46992 225616
rect 57888 225564 57940 225616
rect 56508 225224 56560 225276
rect 57244 225224 57296 225276
rect 381544 224612 381596 224664
rect 384396 224612 384448 224664
rect 51540 223592 51592 223644
rect 55864 223524 55916 223576
rect 52460 223456 52512 223508
rect 56048 223456 56100 223508
rect 57888 222844 57940 222896
rect 65708 222844 65760 222896
rect 57244 222164 57296 222216
rect 60648 222096 60700 222148
rect 44916 220804 44968 220856
rect 47584 220804 47636 220856
rect 56048 220736 56100 220788
rect 56968 220736 57020 220788
rect 65708 220736 65760 220788
rect 69388 220736 69440 220788
rect 394056 220736 394108 220788
rect 396448 220736 396500 220788
rect 368940 220056 368992 220108
rect 377312 220056 377364 220108
rect 77944 218696 77996 218748
rect 87512 218696 87564 218748
rect 69388 218016 69440 218068
rect 118700 218016 118752 218068
rect 580080 218016 580132 218068
rect 71964 217948 72016 218000
rect 45100 217268 45152 217320
rect 53840 217268 53892 217320
rect 380164 216656 380216 216708
rect 381544 216656 381596 216708
rect 45008 216588 45060 216640
rect 46204 216588 46256 216640
rect 56968 216452 57020 216504
rect 59636 216452 59688 216504
rect 71964 215296 72016 215348
rect 76564 215228 76616 215280
rect 53840 214548 53892 214600
rect 77944 214548 77996 214600
rect 358728 214548 358780 214600
rect 368940 214548 368992 214600
rect 3332 213936 3384 213988
rect 179512 213936 179564 213988
rect 60740 213868 60792 213920
rect 63500 213868 63552 213920
rect 59636 213188 59688 213240
rect 68284 213188 68336 213240
rect 47584 212440 47636 212492
rect 52460 212440 52512 212492
rect 55864 212440 55916 212492
rect 59268 212440 59320 212492
rect 344100 211760 344152 211812
rect 358728 211760 358780 211812
rect 63500 211012 63552 211064
rect 65892 211012 65944 211064
rect 87512 209788 87564 209840
rect 95884 209788 95936 209840
rect 159364 209788 159416 209840
rect 162124 209788 162176 209840
rect 392584 209788 392636 209840
rect 394056 209788 394108 209840
rect 59268 209108 59320 209160
rect 62120 209108 62172 209160
rect 46204 208972 46256 209024
rect 48780 208972 48832 209024
rect 68284 208904 68336 208956
rect 75552 208904 75604 208956
rect 52460 208632 52512 208684
rect 55864 208632 55916 208684
rect 65892 208360 65944 208412
rect 376760 208360 376812 208412
rect 380164 208360 380216 208412
rect 71688 208292 71740 208344
rect 341524 207000 341576 207052
rect 344100 207000 344152 207052
rect 389180 207000 389232 207052
rect 392676 207000 392728 207052
rect 62120 205640 62172 205692
rect 48780 205572 48832 205624
rect 56416 205572 56468 205624
rect 189724 205640 189776 205692
rect 580080 205640 580132 205692
rect 66444 205572 66496 205624
rect 76564 205368 76616 205420
rect 78312 205368 78364 205420
rect 377680 204892 377732 204944
rect 389180 204892 389232 204944
rect 71780 204212 71832 204264
rect 73804 204212 73856 204264
rect 56416 202920 56468 202972
rect 62120 202920 62172 202972
rect 374000 202240 374052 202292
rect 377680 202240 377732 202292
rect 147772 202104 147824 202156
rect 176660 202104 176712 202156
rect 3332 201832 3384 201884
rect 7564 201832 7616 201884
rect 62120 201424 62172 201476
rect 64236 201424 64288 201476
rect 66444 201424 66496 201476
rect 69664 201424 69716 201476
rect 75552 201424 75604 201476
rect 76564 201424 76616 201476
rect 77944 201424 77996 201476
rect 80704 201424 80756 201476
rect 78312 201356 78364 201408
rect 79968 201356 80020 201408
rect 375380 201288 375432 201340
rect 376760 201288 376812 201340
rect 155960 199384 156012 199436
rect 296720 199384 296772 199436
rect 351184 199384 351236 199436
rect 374000 199384 374052 199436
rect 338764 198704 338816 198756
rect 341524 198704 341576 198756
rect 73804 198228 73856 198280
rect 75552 198228 75604 198280
rect 148968 197956 149020 198008
rect 207020 197956 207072 198008
rect 154488 197412 154540 197464
rect 155960 197412 156012 197464
rect 79968 197344 80020 197396
rect 84844 197276 84896 197328
rect 152740 197276 152792 197328
rect 157984 197276 158036 197328
rect 138664 196732 138716 196784
rect 164240 196732 164292 196784
rect 151176 196664 151228 196716
rect 236000 196664 236052 196716
rect 155960 196596 156012 196648
rect 327080 196596 327132 196648
rect 162124 196460 162176 196512
rect 164148 196460 164200 196512
rect 367100 196460 367152 196512
rect 375380 196460 375432 196512
rect 56600 195916 56652 195968
rect 138112 195916 138164 195968
rect 160100 195916 160152 195968
rect 386420 195916 386472 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 157616 195848 157668 195900
rect 267004 195848 267056 195900
rect 75552 194624 75604 194676
rect 76656 194624 76708 194676
rect 115940 194556 115992 194608
rect 140780 194556 140832 194608
rect 164148 194488 164200 194540
rect 167644 194488 167696 194540
rect 504456 191836 504508 191888
rect 579804 191836 579856 191888
rect 55864 191768 55916 191820
rect 64144 191768 64196 191820
rect 144460 190476 144512 190528
rect 362224 190476 362276 190528
rect 367008 190476 367060 190528
rect 145012 190272 145064 190324
rect 64236 189728 64288 189780
rect 69756 189728 69808 189780
rect 144644 189048 144696 189100
rect 145012 189048 145064 189100
rect 76564 188164 76616 188216
rect 78588 188164 78640 188216
rect 3332 187688 3384 187740
rect 115204 187688 115256 187740
rect 336004 187688 336056 187740
rect 338764 187688 338816 187740
rect 76656 187348 76708 187400
rect 79968 187348 80020 187400
rect 84844 186940 84896 186992
rect 86224 186940 86276 186992
rect 69664 185988 69716 186040
rect 71044 185988 71096 186040
rect 159548 185852 159600 185904
rect 159916 185512 159968 185564
rect 79968 184832 80020 184884
rect 81440 184832 81492 184884
rect 78680 184764 78732 184816
rect 80796 184764 80848 184816
rect 390560 183472 390612 183524
rect 392584 183472 392636 183524
rect 131764 183404 131816 183456
rect 133972 183404 134024 183456
rect 81440 182180 81492 182232
rect 86316 182112 86368 182164
rect 144644 181092 144696 181144
rect 151912 181024 151964 181076
rect 159916 180684 159968 180736
rect 121460 180140 121512 180192
rect 136364 180140 136416 180192
rect 133972 180072 134024 180124
rect 159916 180072 159968 180124
rect 151912 179460 151964 179512
rect 153936 179460 153988 179512
rect 149060 179392 149112 179444
rect 154396 179392 154448 179444
rect 157800 179392 157852 179444
rect 158628 179392 158680 179444
rect 169760 179392 169812 179444
rect 136732 178780 136784 178832
rect 122840 178644 122892 178696
rect 136456 178644 136508 178696
rect 136364 178372 136416 178424
rect 71044 178304 71096 178356
rect 72424 178304 72476 178356
rect 330024 177964 330076 178016
rect 336004 177964 336056 178016
rect 134984 177760 135036 177812
rect 136640 177760 136692 177812
rect 124220 177284 124272 177336
rect 136456 177284 136508 177336
rect 135260 177216 135312 177268
rect 136548 177216 136600 177268
rect 159916 176400 159968 176452
rect 126980 176128 127032 176180
rect 134984 176128 135036 176180
rect 125600 175992 125652 176044
rect 136364 175992 136416 176044
rect 144092 175992 144144 176044
rect 149336 175992 149388 176044
rect 69756 175924 69808 175976
rect 92480 175924 92532 175976
rect 118884 175924 118936 175976
rect 144460 175788 144512 175840
rect 149980 175788 150032 175840
rect 158168 175720 158220 175772
rect 165068 175924 165120 175976
rect 580080 175924 580132 175976
rect 159180 175856 159232 175908
rect 165160 175856 165212 175908
rect 167000 175856 167052 175908
rect 163504 175720 163556 175772
rect 163596 175652 163648 175704
rect 153936 175380 153988 175432
rect 154396 175380 154448 175432
rect 155500 175244 155552 175296
rect 159180 175380 159232 175432
rect 128360 175176 128412 175228
rect 135260 175176 135312 175228
rect 385684 175176 385736 175228
rect 390468 175176 390520 175228
rect 141608 174768 141660 174820
rect 146484 174768 146536 174820
rect 149060 174768 149112 174820
rect 143080 174700 143132 174752
rect 152372 174700 152424 174752
rect 162492 174700 162544 174752
rect 156512 174632 156564 174684
rect 161480 174564 161532 174616
rect 135904 174360 135956 174412
rect 155500 174496 155552 174548
rect 146484 174292 146536 174344
rect 133880 173884 133932 173936
rect 137376 173884 137428 173936
rect 86316 173816 86368 173868
rect 87972 173816 88024 173868
rect 327724 174088 327776 174140
rect 330024 174088 330076 174140
rect 167644 173816 167696 173868
rect 169116 173816 169168 173868
rect 149336 172932 149388 172984
rect 150440 172932 150492 172984
rect 165436 172932 165488 172984
rect 131120 172524 131172 172576
rect 136548 172524 136600 172576
rect 359832 172456 359884 172508
rect 362224 172456 362276 172508
rect 138020 172116 138072 172168
rect 140780 172116 140832 172168
rect 64144 171776 64196 171828
rect 69940 171776 69992 171828
rect 135260 171640 135312 171692
rect 138664 171640 138716 171692
rect 92480 171368 92532 171420
rect 94504 171368 94556 171420
rect 132500 171096 132552 171148
rect 136732 171096 136784 171148
rect 162860 169940 162912 169992
rect 163504 169940 163556 169992
rect 87972 169804 88024 169856
rect 88984 169804 89036 169856
rect 169116 169736 169168 169788
rect 170404 169736 170456 169788
rect 346308 169736 346360 169788
rect 351184 169736 351236 169788
rect 86224 168852 86276 168904
rect 88340 168852 88392 168904
rect 69940 168240 69992 168292
rect 77208 168240 77260 168292
rect 80704 168240 80756 168292
rect 86868 168240 86920 168292
rect 80796 167016 80848 167068
rect 82084 167016 82136 167068
rect 163596 166336 163648 166388
rect 163596 166132 163648 166184
rect 340144 166064 340196 166116
rect 346308 166064 346360 166116
rect 188344 165588 188396 165640
rect 580080 165588 580132 165640
rect 88340 165520 88392 165572
rect 90364 165520 90416 165572
rect 356704 165316 356756 165368
rect 359832 165316 359884 165368
rect 77208 164840 77260 164892
rect 85212 164840 85264 164892
rect 118976 164840 119028 164892
rect 580816 164840 580868 164892
rect 86868 164160 86920 164212
rect 91560 164160 91612 164212
rect 155224 164160 155276 164212
rect 160100 164160 160152 164212
rect 3332 162868 3384 162920
rect 181260 162868 181312 162920
rect 85212 162800 85264 162852
rect 91744 162800 91796 162852
rect 20076 162120 20128 162172
rect 182916 162120 182968 162172
rect 324320 161440 324372 161492
rect 327724 161440 327776 161492
rect 170404 160692 170456 160744
rect 173900 160692 173952 160744
rect 72424 160420 72476 160472
rect 76748 160420 76800 160472
rect 94504 160080 94556 160132
rect 163688 160080 163740 160132
rect 166264 160080 166316 160132
rect 382280 160080 382332 160132
rect 385684 160080 385736 160132
rect 98644 160012 98696 160064
rect 91560 159332 91612 159384
rect 98184 159332 98236 159384
rect 319904 158720 319956 158772
rect 324320 158720 324372 158772
rect 82084 158040 82136 158092
rect 83464 158040 83516 158092
rect 160100 158040 160152 158092
rect 166356 158040 166408 158092
rect 119068 157972 119120 158024
rect 580172 157972 580224 158024
rect 173900 157632 173952 157684
rect 175924 157632 175976 157684
rect 76748 155864 76800 155916
rect 79324 155864 79376 155916
rect 353944 155864 353996 155916
rect 356704 155932 356756 155984
rect 374644 155864 374696 155916
rect 382188 155932 382240 155984
rect 303988 155184 304040 155236
rect 319904 155184 319956 155236
rect 322204 155184 322256 155236
rect 340144 155184 340196 155236
rect 98184 153144 98236 153196
rect 102784 153144 102836 153196
rect 301504 152804 301556 152856
rect 303988 152804 304040 152856
rect 180064 151784 180116 151836
rect 579988 151784 580040 151836
rect 88984 150424 89036 150476
rect 372620 150424 372672 150476
rect 374644 150424 374696 150476
rect 94780 150356 94832 150408
rect 3240 149676 3292 149728
rect 22928 149676 22980 149728
rect 91744 148316 91796 148368
rect 109684 148316 109736 148368
rect 134064 147636 134116 147688
rect 135904 147636 135956 147688
rect 45560 146956 45612 147008
rect 48964 146956 49016 147008
rect 166356 146956 166408 147008
rect 168380 146956 168432 147008
rect 166264 146888 166316 146940
rect 180156 146888 180208 146940
rect 94780 146276 94832 146328
rect 371884 146276 371936 146328
rect 372620 146276 372672 146328
rect 97264 146208 97316 146260
rect 141700 146208 141752 146260
rect 142436 146208 142488 146260
rect 350540 144780 350592 144832
rect 353944 144780 353996 144832
rect 33784 144440 33836 144492
rect 182640 144440 182692 144492
rect 10416 144372 10468 144424
rect 182548 144372 182600 144424
rect 6184 144304 6236 144356
rect 182272 144304 182324 144356
rect 118332 144236 118384 144288
rect 398196 144236 398248 144288
rect 118240 144168 118292 144220
rect 398104 144168 398156 144220
rect 98644 143488 98696 143540
rect 100944 143488 100996 143540
rect 146484 143488 146536 143540
rect 148048 143488 148100 143540
rect 153476 143488 153528 143540
rect 158996 143488 159048 143540
rect 147680 143420 147732 143472
rect 149612 143420 149664 143472
rect 152464 143420 152516 143472
rect 157432 143420 157484 143472
rect 137744 143352 137796 143404
rect 139584 143352 139636 143404
rect 163596 143148 163648 143200
rect 174636 143148 174688 143200
rect 150532 143080 150584 143132
rect 154580 143080 154632 143132
rect 164516 143080 164568 143132
rect 176200 143080 176252 143132
rect 122840 143012 122892 143064
rect 134064 143012 134116 143064
rect 144460 143012 144512 143064
rect 160560 143012 160612 143064
rect 163504 143012 163556 143064
rect 178040 143012 178092 143064
rect 118516 142944 118568 142996
rect 398380 142944 398432 142996
rect 118424 142876 118476 142928
rect 398288 142876 398340 142928
rect 102784 142808 102836 142860
rect 108304 142808 108356 142860
rect 120724 142808 120776 142860
rect 477500 142808 477552 142860
rect 140688 142128 140740 142180
rect 142160 142128 142212 142180
rect 149520 142128 149572 142180
rect 152740 142128 152792 142180
rect 157340 142128 157392 142180
rect 163688 142128 163740 142180
rect 175924 142128 175976 142180
rect 181168 142060 181220 142112
rect 40040 141652 40092 141704
rect 180984 141652 181036 141704
rect 4896 141584 4948 141636
rect 182456 141584 182508 141636
rect 118148 141516 118200 141568
rect 542360 141516 542412 141568
rect 119252 141448 119304 141500
rect 580264 141448 580316 141500
rect 119160 141380 119212 141432
rect 580540 141380 580592 141432
rect 121276 140428 121328 140480
rect 122840 140428 122892 140480
rect 79324 140292 79376 140344
rect 82728 140292 82780 140344
rect 100944 140292 100996 140344
rect 181076 140292 181128 140344
rect 10324 140224 10376 140276
rect 182732 140224 182784 140276
rect 4804 140156 4856 140208
rect 182364 140156 182416 140208
rect 83464 140088 83516 140140
rect 85028 140088 85080 140140
rect 119988 140088 120040 140140
rect 301504 140088 301556 140140
rect 118056 140020 118108 140072
rect 412640 140020 412692 140072
rect 90364 139816 90416 139868
rect 91468 139816 91520 139868
rect 118608 139476 118660 139528
rect 178224 139476 178276 139528
rect 43444 139408 43496 139460
rect 182180 139408 182232 139460
rect 369768 139408 369820 139460
rect 371884 139408 371936 139460
rect 178224 139340 178276 139392
rect 580172 139340 580224 139392
rect 4068 138660 4120 138712
rect 25504 138660 25556 138712
rect 85028 138048 85080 138100
rect 86224 138048 86276 138100
rect 367744 137980 367796 138032
rect 369768 137980 369820 138032
rect 4068 136688 4120 136740
rect 117320 136688 117372 136740
rect 3332 136620 3384 136672
rect 119344 136620 119396 136672
rect 345664 136552 345716 136604
rect 350540 136620 350592 136672
rect 117964 136144 118016 136196
rect 119988 136144 120040 136196
rect 3332 135260 3384 135312
rect 117320 135260 117372 135312
rect 91468 135192 91520 135244
rect 93768 135192 93820 135244
rect 82820 134852 82872 134904
rect 85212 134852 85264 134904
rect 295984 134512 296036 134564
rect 322204 134512 322256 134564
rect 3240 133900 3292 133952
rect 117320 133900 117372 133952
rect 108304 133152 108356 133204
rect 117780 133152 117832 133204
rect 25504 132404 25556 132456
rect 117320 132404 117372 132456
rect 86224 131112 86276 131164
rect 89536 131112 89588 131164
rect 180156 131112 180208 131164
rect 182180 131112 182232 131164
rect 365720 131112 365772 131164
rect 367744 131112 367796 131164
rect 7564 131044 7616 131096
rect 117320 131044 117372 131096
rect 93860 130092 93912 130144
rect 95608 130092 95660 130144
rect 22836 129684 22888 129736
rect 117320 129684 117372 129736
rect 89536 129616 89588 129668
rect 92388 129616 92440 129668
rect 97264 128596 97316 128648
rect 99748 128596 99800 128648
rect 109684 128324 109736 128376
rect 112444 128324 112496 128376
rect 22928 128256 22980 128308
rect 117320 128256 117372 128308
rect 363604 127712 363656 127764
rect 365720 127712 365772 127764
rect 22744 126896 22796 126948
rect 117320 126896 117372 126948
rect 85212 126828 85264 126880
rect 88800 126828 88852 126880
rect 182824 125604 182876 125656
rect 580172 125604 580224 125656
rect 8944 125536 8996 125588
rect 117320 125536 117372 125588
rect 95608 125468 95660 125520
rect 97172 125468 97224 125520
rect 4988 124108 5040 124160
rect 117320 124108 117372 124160
rect 342260 124108 342312 124160
rect 345664 124176 345716 124228
rect 88800 124040 88852 124092
rect 92388 124040 92440 124092
rect 99748 124040 99800 124092
rect 102048 124040 102100 124092
rect 92480 123428 92532 123480
rect 100760 123428 100812 123480
rect 24124 122748 24176 122800
rect 117320 122748 117372 122800
rect 100760 121796 100812 121848
rect 102140 121796 102192 121848
rect 92388 121728 92440 121780
rect 94412 121728 94464 121780
rect 37924 121388 37976 121440
rect 117320 121388 117372 121440
rect 97172 120844 97224 120896
rect 105728 120844 105780 120896
rect 19984 120028 20036 120080
rect 117320 120028 117372 120080
rect 102048 119960 102100 120012
rect 104348 119960 104400 120012
rect 15844 118600 15896 118652
rect 117320 118600 117372 118652
rect 117964 118600 118016 118652
rect 102140 118532 102192 118584
rect 104716 118532 104768 118584
rect 112444 118532 112496 118584
rect 115480 118532 115532 118584
rect 104348 118396 104400 118448
rect 108304 118396 108356 118448
rect 118056 118396 118108 118448
rect 94412 118260 94464 118312
rect 97172 118260 97224 118312
rect 48964 117920 49016 117972
rect 63500 117920 63552 117972
rect 360200 117648 360252 117700
rect 363604 117648 363656 117700
rect 23480 117240 23532 117292
rect 117320 117240 117372 117292
rect 293224 116968 293276 117020
rect 295984 116968 296036 117020
rect 97172 115948 97224 116000
rect 95884 115880 95936 115932
rect 98644 115880 98696 115932
rect 100668 115880 100720 115932
rect 105728 115880 105780 115932
rect 110328 115880 110380 115932
rect 115480 115880 115532 115932
rect 117780 115880 117832 115932
rect 338764 115880 338816 115932
rect 342260 115948 342312 116000
rect 358268 115064 358320 115116
rect 360200 115064 360252 115116
rect 63500 114452 63552 114504
rect 117320 114452 117372 114504
rect 117688 114452 117740 114504
rect 120908 114452 120960 114504
rect 104716 114384 104768 114436
rect 107936 114384 107988 114436
rect 351920 113772 351972 113824
rect 358268 113772 358320 113824
rect 110328 113092 110380 113144
rect 117320 113092 117372 113144
rect 336740 111868 336792 111920
rect 338764 111868 338816 111920
rect 349160 111868 349212 111920
rect 351920 111868 351972 111920
rect 180156 111800 180208 111852
rect 580172 111800 580224 111852
rect 3148 111732 3200 111784
rect 43444 111732 43496 111784
rect 100668 111732 100720 111784
rect 117320 111732 117372 111784
rect 183284 111732 183336 111784
rect 336740 111732 336792 111784
rect 107936 110440 107988 110492
rect 117320 110372 117372 110424
rect 183468 110372 183520 110424
rect 349160 110440 349212 110492
rect 183376 108944 183428 108996
rect 410524 108944 410576 108996
rect 183468 106224 183520 106276
rect 409144 106224 409196 106276
rect 183468 104796 183520 104848
rect 407764 104796 407816 104848
rect 183468 103436 183520 103488
rect 406384 103436 406436 103488
rect 183468 102076 183520 102128
rect 405004 102076 405056 102128
rect 98644 100648 98696 100700
rect 100760 100648 100812 100700
rect 183468 100648 183520 100700
rect 403624 100648 403676 100700
rect 183468 99288 183520 99340
rect 400864 99288 400916 99340
rect 108304 98676 108356 98728
rect 109684 98676 109736 98728
rect 117780 97928 117832 97980
rect 120908 97928 120960 97980
rect 183468 97928 183520 97980
rect 399484 97928 399536 97980
rect 100760 97248 100812 97300
rect 109776 97248 109828 97300
rect 183192 96568 183244 96620
rect 418804 96568 418856 96620
rect 183284 95140 183336 95192
rect 417424 95140 417476 95192
rect 183284 93780 183336 93832
rect 414664 93780 414716 93832
rect 109776 93576 109828 93628
rect 113824 93576 113876 93628
rect 109684 93236 109736 93288
rect 110420 93236 110472 93288
rect 183468 92420 183520 92472
rect 413284 92420 413336 92472
rect 110420 91060 110472 91112
rect 115296 90992 115348 91044
rect 183468 89632 183520 89684
rect 189724 89632 189776 89684
rect 183468 88204 183520 88256
rect 188344 88204 188396 88256
rect 3148 85552 3200 85604
rect 3516 85552 3568 85604
rect 3608 85552 3660 85604
rect 183468 85552 183520 85604
rect 580172 85552 580224 85604
rect 3608 85348 3660 85400
rect 3884 84940 3936 84992
rect 3056 84804 3108 84856
rect 3332 84804 3384 84856
rect 3884 84668 3936 84720
rect 3976 84192 4028 84244
rect 120448 84192 120500 84244
rect 178960 82084 179012 82136
rect 580356 82084 580408 82136
rect 183468 81404 183520 81456
rect 555424 81404 555476 81456
rect 113824 80656 113876 80708
rect 119344 79976 119396 80028
rect 125048 80248 125100 80300
rect 123668 80044 123720 80096
rect 124956 79908 125008 79960
rect 122932 79840 122984 79892
rect 126014 79840 126066 79892
rect 126290 79840 126342 79892
rect 125508 79772 125560 79824
rect 125922 79772 125974 79824
rect 126060 79704 126112 79756
rect 126336 79704 126388 79756
rect 126750 79908 126802 79960
rect 126566 79840 126618 79892
rect 126658 79840 126710 79892
rect 126934 79908 126986 79960
rect 127026 79908 127078 79960
rect 127486 79908 127538 79960
rect 127762 79908 127814 79960
rect 128038 79908 128090 79960
rect 128222 79908 128274 79960
rect 128406 79908 128458 79960
rect 5172 79568 5224 79620
rect 120724 79568 120776 79620
rect 115204 79432 115256 79484
rect 125876 79500 125928 79552
rect 125968 79500 126020 79552
rect 127072 79772 127124 79824
rect 126980 79704 127032 79756
rect 127670 79840 127722 79892
rect 126888 79636 126940 79688
rect 127164 79500 127216 79552
rect 128084 79772 128136 79824
rect 128176 79772 128228 79824
rect 128360 79568 128412 79620
rect 129050 79908 129102 79960
rect 129142 79908 129194 79960
rect 129326 79908 129378 79960
rect 129602 79908 129654 79960
rect 129694 79908 129746 79960
rect 129786 79908 129838 79960
rect 129970 79908 130022 79960
rect 128958 79840 129010 79892
rect 129418 79840 129470 79892
rect 129510 79840 129562 79892
rect 128912 79704 128964 79756
rect 129096 79704 129148 79756
rect 129280 79636 129332 79688
rect 129372 79636 129424 79688
rect 130154 79840 130206 79892
rect 130246 79840 130298 79892
rect 129786 79772 129838 79824
rect 129832 79636 129884 79688
rect 129924 79636 129976 79688
rect 130200 79704 130252 79756
rect 130522 79908 130574 79960
rect 129464 79568 129516 79620
rect 129556 79568 129608 79620
rect 130016 79568 130068 79620
rect 130476 79636 130528 79688
rect 128544 79500 128596 79552
rect 130982 79908 131034 79960
rect 131534 79908 131586 79960
rect 131718 79908 131770 79960
rect 130890 79840 130942 79892
rect 130936 79704 130988 79756
rect 131166 79840 131218 79892
rect 131350 79840 131402 79892
rect 131212 79636 131264 79688
rect 131488 79772 131540 79824
rect 131994 79840 132046 79892
rect 132270 79840 132322 79892
rect 132454 79840 132506 79892
rect 131810 79772 131862 79824
rect 131672 79704 131724 79756
rect 131764 79636 131816 79688
rect 131028 79500 131080 79552
rect 132040 79500 132092 79552
rect 132546 79772 132598 79824
rect 132408 79636 132460 79688
rect 132914 79908 132966 79960
rect 133926 79908 133978 79960
rect 134110 79908 134162 79960
rect 134294 79908 134346 79960
rect 135030 79908 135082 79960
rect 135122 79908 135174 79960
rect 135490 79908 135542 79960
rect 132822 79840 132874 79892
rect 133190 79840 133242 79892
rect 133742 79840 133794 79892
rect 132592 79568 132644 79620
rect 132684 79500 132736 79552
rect 132776 79500 132828 79552
rect 133052 79500 133104 79552
rect 133374 79772 133426 79824
rect 133650 79772 133702 79824
rect 133604 79568 133656 79620
rect 133880 79772 133932 79824
rect 134064 79636 134116 79688
rect 134156 79568 134208 79620
rect 134570 79840 134622 79892
rect 134754 79840 134806 79892
rect 134432 79568 134484 79620
rect 133328 79500 133380 79552
rect 133696 79500 133748 79552
rect 133972 79500 134024 79552
rect 134984 79568 135036 79620
rect 135076 79568 135128 79620
rect 134064 79432 134116 79484
rect 120724 79364 120776 79416
rect 125324 79296 125376 79348
rect 126244 79296 126296 79348
rect 134524 79296 134576 79348
rect 135306 79772 135358 79824
rect 135674 79840 135726 79892
rect 135628 79636 135680 79688
rect 136594 79908 136646 79960
rect 137422 79908 137474 79960
rect 137514 79908 137566 79960
rect 137606 79908 137658 79960
rect 137698 79908 137750 79960
rect 138066 79908 138118 79960
rect 138526 79908 138578 79960
rect 138618 79908 138670 79960
rect 136134 79840 136186 79892
rect 136318 79840 136370 79892
rect 136410 79840 136462 79892
rect 136962 79840 137014 79892
rect 137054 79840 137106 79892
rect 137238 79840 137290 79892
rect 135536 79500 135588 79552
rect 135996 79500 136048 79552
rect 135352 79364 135404 79416
rect 136502 79772 136554 79824
rect 136778 79772 136830 79824
rect 136870 79772 136922 79824
rect 136732 79636 136784 79688
rect 136548 79568 136600 79620
rect 136272 79500 136324 79552
rect 136364 79500 136416 79552
rect 137100 79704 137152 79756
rect 137284 79704 137336 79756
rect 137376 79636 137428 79688
rect 136916 79568 136968 79620
rect 137008 79500 137060 79552
rect 137468 79500 137520 79552
rect 136732 79432 136784 79484
rect 138158 79840 138210 79892
rect 138250 79840 138302 79892
rect 138020 79636 138072 79688
rect 139262 79908 139314 79960
rect 139354 79908 139406 79960
rect 139446 79908 139498 79960
rect 138480 79568 138532 79620
rect 138388 79500 138440 79552
rect 138894 79840 138946 79892
rect 138756 79568 138808 79620
rect 139078 79772 139130 79824
rect 139032 79568 139084 79620
rect 139124 79568 139176 79620
rect 138940 79432 138992 79484
rect 139446 79772 139498 79824
rect 139814 79908 139866 79960
rect 140090 79908 140142 79960
rect 140274 79908 140326 79960
rect 140366 79908 140418 79960
rect 140550 79908 140602 79960
rect 140734 79908 140786 79960
rect 140826 79908 140878 79960
rect 141194 79908 141246 79960
rect 141286 79908 141338 79960
rect 141378 79908 141430 79960
rect 141562 79908 141614 79960
rect 141654 79908 141706 79960
rect 139630 79840 139682 79892
rect 139906 79840 139958 79892
rect 139492 79636 139544 79688
rect 139860 79704 139912 79756
rect 139952 79704 140004 79756
rect 140320 79772 140372 79824
rect 140918 79840 140970 79892
rect 141010 79840 141062 79892
rect 140688 79704 140740 79756
rect 140780 79704 140832 79756
rect 140596 79636 140648 79688
rect 140228 79568 140280 79620
rect 140872 79568 140924 79620
rect 141056 79568 141108 79620
rect 139768 79500 139820 79552
rect 140964 79500 141016 79552
rect 141470 79840 141522 79892
rect 139952 79432 140004 79484
rect 141608 79568 141660 79620
rect 141930 79908 141982 79960
rect 141516 79500 141568 79552
rect 141700 79500 141752 79552
rect 142206 79908 142258 79960
rect 142390 79908 142442 79960
rect 142482 79908 142534 79960
rect 142574 79908 142626 79960
rect 142666 79908 142718 79960
rect 143218 79908 143270 79960
rect 142712 79772 142764 79824
rect 142942 79772 142994 79824
rect 143034 79772 143086 79824
rect 143126 79772 143178 79824
rect 142804 79636 142856 79688
rect 142252 79568 142304 79620
rect 142068 79500 142120 79552
rect 142988 79636 143040 79688
rect 143172 79636 143224 79688
rect 143264 79636 143316 79688
rect 143080 79568 143132 79620
rect 143770 79908 143822 79960
rect 143862 79908 143914 79960
rect 144138 79840 144190 79892
rect 144046 79772 144098 79824
rect 144414 79908 144466 79960
rect 144506 79908 144558 79960
rect 144690 79908 144742 79960
rect 143908 79568 143960 79620
rect 144092 79568 144144 79620
rect 144184 79568 144236 79620
rect 144276 79568 144328 79620
rect 143448 79500 143500 79552
rect 143540 79500 143592 79552
rect 144552 79704 144604 79756
rect 144644 79704 144696 79756
rect 144966 79772 145018 79824
rect 145150 79908 145202 79960
rect 145426 79908 145478 79960
rect 145794 79908 145846 79960
rect 145886 79908 145938 79960
rect 144920 79636 144972 79688
rect 145012 79636 145064 79688
rect 144828 79568 144880 79620
rect 145610 79840 145662 79892
rect 145840 79772 145892 79824
rect 145656 79636 145708 79688
rect 147082 79908 147134 79960
rect 147450 79908 147502 79960
rect 148094 79908 148146 79960
rect 148186 79908 148238 79960
rect 148278 79908 148330 79960
rect 149014 79908 149066 79960
rect 149106 79908 149158 79960
rect 146990 79840 147042 79892
rect 146622 79772 146674 79824
rect 147266 79840 147318 79892
rect 147910 79840 147962 79892
rect 147404 79772 147456 79824
rect 147726 79772 147778 79824
rect 147818 79772 147870 79824
rect 147128 79636 147180 79688
rect 147220 79568 147272 79620
rect 147956 79704 148008 79756
rect 148048 79704 148100 79756
rect 147864 79636 147916 79688
rect 147772 79568 147824 79620
rect 145380 79500 145432 79552
rect 146024 79500 146076 79552
rect 146300 79500 146352 79552
rect 147496 79500 147548 79552
rect 148370 79840 148422 79892
rect 148830 79840 148882 79892
rect 148278 79772 148330 79824
rect 148784 79704 148836 79756
rect 148324 79636 148376 79688
rect 149474 79908 149526 79960
rect 149750 79908 149802 79960
rect 149382 79840 149434 79892
rect 149060 79636 149112 79688
rect 149244 79636 149296 79688
rect 149796 79636 149848 79688
rect 150026 79908 150078 79960
rect 148876 79568 148928 79620
rect 149520 79500 149572 79552
rect 149888 79568 149940 79620
rect 150118 79840 150170 79892
rect 150164 79704 150216 79756
rect 150486 79908 150538 79960
rect 150762 79908 150814 79960
rect 151222 79908 151274 79960
rect 151498 79908 151550 79960
rect 151590 79908 151642 79960
rect 151682 79908 151734 79960
rect 150348 79568 150400 79620
rect 150946 79772 150998 79824
rect 150808 79636 150860 79688
rect 150900 79636 150952 79688
rect 150992 79636 151044 79688
rect 151176 79568 151228 79620
rect 151958 79908 152010 79960
rect 152050 79908 152102 79960
rect 152142 79908 152194 79960
rect 152510 79908 152562 79960
rect 152970 79908 153022 79960
rect 151866 79840 151918 79892
rect 151820 79704 151872 79756
rect 151912 79568 151964 79620
rect 151544 79500 151596 79552
rect 151728 79500 151780 79552
rect 152694 79840 152746 79892
rect 152556 79772 152608 79824
rect 152464 79568 152516 79620
rect 178500 80724 178552 80776
rect 393964 80724 394016 80776
rect 174728 80656 174780 80708
rect 174544 80520 174596 80572
rect 176016 80520 176068 80572
rect 504456 80656 504508 80708
rect 176108 80452 176160 80504
rect 175280 80384 175332 80436
rect 182180 80384 182232 80436
rect 153246 79908 153298 79960
rect 153016 79636 153068 79688
rect 152924 79568 152976 79620
rect 152740 79500 152792 79552
rect 144000 79432 144052 79484
rect 151452 79432 151504 79484
rect 153614 79908 153666 79960
rect 153798 79908 153850 79960
rect 153706 79840 153758 79892
rect 153522 79772 153574 79824
rect 153660 79704 153712 79756
rect 153568 79636 153620 79688
rect 153292 79568 153344 79620
rect 154074 79908 154126 79960
rect 154166 79772 154218 79824
rect 153936 79636 153988 79688
rect 154120 79636 154172 79688
rect 153844 79500 153896 79552
rect 154212 79500 154264 79552
rect 154626 79908 154678 79960
rect 154994 79908 155046 79960
rect 155178 79908 155230 79960
rect 155270 79908 155322 79960
rect 156006 79908 156058 79960
rect 156282 79908 156334 79960
rect 154718 79840 154770 79892
rect 154580 79636 154632 79688
rect 154948 79772 155000 79824
rect 155454 79840 155506 79892
rect 155822 79840 155874 79892
rect 155914 79840 155966 79892
rect 155224 79636 155276 79688
rect 155316 79636 155368 79688
rect 155408 79636 155460 79688
rect 154764 79568 154816 79620
rect 156190 79840 156242 79892
rect 156006 79772 156058 79824
rect 156144 79636 156196 79688
rect 156236 79568 156288 79620
rect 156466 79908 156518 79960
rect 157202 79908 157254 79960
rect 157754 79908 157806 79960
rect 157846 79908 157898 79960
rect 158030 79908 158082 79960
rect 155132 79432 155184 79484
rect 155776 79432 155828 79484
rect 140504 79364 140556 79416
rect 141332 79364 141384 79416
rect 141424 79364 141476 79416
rect 141884 79364 141936 79416
rect 142068 79364 142120 79416
rect 146944 79364 146996 79416
rect 149704 79364 149756 79416
rect 156328 79500 156380 79552
rect 156558 79840 156610 79892
rect 157018 79840 157070 79892
rect 156834 79772 156886 79824
rect 156926 79772 156978 79824
rect 157156 79772 157208 79824
rect 156512 79704 156564 79756
rect 156604 79704 156656 79756
rect 156880 79636 156932 79688
rect 157064 79568 157116 79620
rect 157386 79840 157438 79892
rect 157662 79840 157714 79892
rect 157340 79568 157392 79620
rect 157708 79568 157760 79620
rect 157524 79500 157576 79552
rect 158214 79908 158266 79960
rect 158306 79908 158358 79960
rect 158490 79908 158542 79960
rect 157892 79568 157944 79620
rect 158076 79568 158128 79620
rect 158444 79704 158496 79756
rect 158766 79908 158818 79960
rect 158858 79908 158910 79960
rect 159042 79908 159094 79960
rect 158536 79636 158588 79688
rect 158858 79772 158910 79824
rect 159226 79908 159278 79960
rect 159318 79908 159370 79960
rect 159502 79908 159554 79960
rect 159594 79908 159646 79960
rect 159088 79636 159140 79688
rect 159410 79840 159462 79892
rect 159364 79636 159416 79688
rect 159180 79568 159232 79620
rect 159272 79568 159324 79620
rect 158168 79500 158220 79552
rect 158904 79500 158956 79552
rect 159686 79840 159738 79892
rect 159962 79840 160014 79892
rect 160146 79840 160198 79892
rect 159732 79704 159784 79756
rect 160008 79636 160060 79688
rect 156420 79432 156472 79484
rect 138296 79296 138348 79348
rect 146944 79160 146996 79212
rect 149704 79160 149756 79212
rect 153752 79296 153804 79348
rect 153936 79296 153988 79348
rect 154856 79296 154908 79348
rect 155132 79296 155184 79348
rect 156972 79364 157024 79416
rect 157616 79364 157668 79416
rect 159916 79364 159968 79416
rect 160330 79908 160382 79960
rect 160422 79908 160474 79960
rect 160698 79908 160750 79960
rect 161066 79908 161118 79960
rect 161158 79908 161210 79960
rect 161250 79908 161302 79960
rect 160606 79840 160658 79892
rect 160468 79772 160520 79824
rect 160376 79704 160428 79756
rect 160284 79568 160336 79620
rect 160560 79636 160612 79688
rect 160652 79568 160704 79620
rect 160974 79840 161026 79892
rect 161020 79704 161072 79756
rect 161112 79704 161164 79756
rect 161204 79636 161256 79688
rect 161802 79908 161854 79960
rect 161894 79908 161946 79960
rect 161618 79840 161670 79892
rect 161434 79772 161486 79824
rect 161572 79704 161624 79756
rect 162078 79908 162130 79960
rect 161940 79772 161992 79824
rect 162262 79840 162314 79892
rect 162354 79840 162406 79892
rect 162446 79840 162498 79892
rect 161848 79704 161900 79756
rect 162032 79704 162084 79756
rect 161480 79636 161532 79688
rect 161756 79636 161808 79688
rect 162308 79636 162360 79688
rect 161296 79568 161348 79620
rect 162124 79568 162176 79620
rect 162906 79840 162958 79892
rect 163274 79840 163326 79892
rect 163228 79704 163280 79756
rect 174452 80316 174504 80368
rect 180156 80316 180208 80368
rect 162676 79636 162728 79688
rect 162768 79636 162820 79688
rect 163320 79636 163372 79688
rect 163412 79636 163464 79688
rect 162492 79568 162544 79620
rect 163918 79908 163970 79960
rect 164194 79908 164246 79960
rect 164838 79908 164890 79960
rect 164930 79908 164982 79960
rect 163642 79840 163694 79892
rect 163734 79840 163786 79892
rect 160836 79500 160888 79552
rect 161664 79500 161716 79552
rect 162400 79500 162452 79552
rect 163136 79500 163188 79552
rect 163412 79500 163464 79552
rect 163964 79772 164016 79824
rect 163780 79704 163832 79756
rect 164148 79636 164200 79688
rect 164700 79568 164752 79620
rect 164884 79568 164936 79620
rect 163964 79500 164016 79552
rect 164332 79500 164384 79552
rect 165758 79908 165810 79960
rect 165850 79908 165902 79960
rect 166034 79908 166086 79960
rect 166310 79908 166362 79960
rect 167414 79908 167466 79960
rect 165942 79840 165994 79892
rect 165804 79704 165856 79756
rect 166034 79772 166086 79824
rect 166126 79772 166178 79824
rect 165896 79636 165948 79688
rect 165712 79568 165764 79620
rect 166954 79840 167006 79892
rect 167138 79840 167190 79892
rect 166172 79636 166224 79688
rect 166356 79636 166408 79688
rect 167368 79772 167420 79824
rect 167184 79636 167236 79688
rect 168058 79908 168110 79960
rect 168334 79908 168386 79960
rect 168150 79840 168202 79892
rect 168518 79840 168570 79892
rect 168610 79840 168662 79892
rect 168702 79840 168754 79892
rect 168380 79704 168432 79756
rect 168472 79704 168524 79756
rect 169530 79908 169582 79960
rect 169990 79840 170042 79892
rect 170358 79840 170410 79892
rect 170818 79840 170870 79892
rect 174636 80248 174688 80300
rect 200120 80248 200172 80300
rect 174452 80180 174504 80232
rect 174544 80180 174596 80232
rect 231860 80180 231912 80232
rect 176016 80112 176068 80164
rect 176108 80112 176160 80164
rect 252560 80112 252612 80164
rect 171094 79908 171146 79960
rect 171278 79908 171330 79960
rect 170726 79772 170778 79824
rect 171554 79840 171606 79892
rect 171738 79840 171790 79892
rect 171232 79772 171284 79824
rect 171370 79772 171422 79824
rect 170864 79704 170916 79756
rect 171508 79704 171560 79756
rect 168104 79636 168156 79688
rect 168196 79636 168248 79688
rect 168656 79636 168708 79688
rect 169024 79636 169076 79688
rect 169484 79636 169536 79688
rect 169944 79636 169996 79688
rect 170634 79636 170686 79688
rect 171140 79636 171192 79688
rect 171600 79636 171652 79688
rect 166080 79568 166132 79620
rect 166632 79568 166684 79620
rect 166908 79568 166960 79620
rect 172382 79908 172434 79960
rect 172566 79840 172618 79892
rect 172658 79840 172710 79892
rect 172934 79840 172986 79892
rect 172336 79772 172388 79824
rect 172520 79704 172572 79756
rect 166540 79500 166592 79552
rect 172244 79568 172296 79620
rect 168748 79500 168800 79552
rect 171508 79500 171560 79552
rect 161848 79432 161900 79484
rect 164516 79432 164568 79484
rect 164700 79432 164752 79484
rect 165068 79432 165120 79484
rect 172428 79432 172480 79484
rect 172612 79568 172664 79620
rect 172704 79432 172756 79484
rect 174544 79976 174596 80028
rect 175188 80044 175240 80096
rect 430580 80044 430632 80096
rect 178408 79976 178460 80028
rect 173578 79908 173630 79960
rect 173670 79908 173722 79960
rect 173946 79908 173998 79960
rect 173210 79840 173262 79892
rect 173670 79772 173722 79824
rect 173256 79704 173308 79756
rect 174130 79840 174182 79892
rect 174176 79704 174228 79756
rect 173624 79636 173676 79688
rect 173808 79568 173860 79620
rect 174728 79432 174780 79484
rect 171784 79364 171836 79416
rect 172152 79364 172204 79416
rect 175280 79364 175332 79416
rect 159640 79296 159692 79348
rect 161940 79296 161992 79348
rect 163412 79296 163464 79348
rect 150348 79228 150400 79280
rect 164516 79228 164568 79280
rect 165068 79228 165120 79280
rect 166632 79296 166684 79348
rect 167000 79296 167052 79348
rect 167460 79296 167512 79348
rect 178040 79364 178092 79416
rect 179420 79296 179472 79348
rect 580448 79296 580500 79348
rect 174176 79228 174228 79280
rect 120448 79092 120500 79144
rect 5080 78820 5132 78872
rect 150348 79092 150400 79144
rect 151452 79092 151504 79144
rect 161848 79092 161900 79144
rect 145196 79024 145248 79076
rect 147588 79024 147640 79076
rect 148968 79024 149020 79076
rect 157248 78956 157300 79008
rect 160560 79024 160612 79076
rect 161296 79024 161348 79076
rect 163504 79092 163556 79144
rect 174268 79160 174320 79212
rect 166540 79092 166592 79144
rect 166908 79092 166960 79144
rect 195980 79092 196032 79144
rect 165068 79024 165120 79076
rect 249800 79024 249852 79076
rect 164516 78956 164568 79008
rect 165620 78956 165672 79008
rect 144460 78888 144512 78940
rect 146944 78888 146996 78940
rect 155040 78888 155092 78940
rect 155500 78888 155552 78940
rect 157708 78888 157760 78940
rect 157984 78888 158036 78940
rect 159364 78888 159416 78940
rect 160284 78888 160336 78940
rect 161664 78888 161716 78940
rect 162216 78888 162268 78940
rect 162584 78888 162636 78940
rect 162952 78888 163004 78940
rect 164240 78888 164292 78940
rect 164792 78888 164844 78940
rect 165712 78888 165764 78940
rect 166080 78888 166132 78940
rect 166540 78956 166592 79008
rect 167000 78956 167052 79008
rect 171324 78956 171376 79008
rect 171692 78956 171744 79008
rect 213920 78956 213972 79008
rect 134064 78820 134116 78872
rect 144000 78820 144052 78872
rect 145196 78820 145248 78872
rect 145656 78820 145708 78872
rect 148324 78820 148376 78872
rect 148508 78820 148560 78872
rect 159180 78820 159232 78872
rect 166632 78820 166684 78872
rect 157616 78752 157668 78804
rect 158076 78752 158128 78804
rect 160192 78752 160244 78804
rect 160928 78752 160980 78804
rect 161572 78752 161624 78804
rect 161940 78752 161992 78804
rect 162216 78752 162268 78804
rect 165068 78752 165120 78804
rect 165804 78752 165856 78804
rect 166080 78752 166132 78804
rect 267740 78888 267792 78940
rect 167000 78820 167052 78872
rect 171876 78820 171928 78872
rect 172520 78820 172572 78872
rect 293224 78820 293276 78872
rect 168288 78752 168340 78804
rect 170496 78752 170548 78804
rect 170864 78752 170916 78804
rect 171784 78752 171836 78804
rect 444380 78752 444432 78804
rect 115296 78684 115348 78736
rect 131580 78684 131632 78736
rect 133880 78684 133932 78736
rect 146852 78684 146904 78736
rect 147312 78684 147364 78736
rect 147956 78684 148008 78736
rect 148140 78684 148192 78736
rect 148324 78684 148376 78736
rect 148692 78684 148744 78736
rect 119988 78616 120040 78668
rect 145656 78616 145708 78668
rect 146024 78616 146076 78668
rect 146392 78616 146444 78668
rect 146760 78616 146812 78668
rect 147588 78616 147640 78668
rect 159180 78684 159232 78736
rect 161848 78684 161900 78736
rect 162124 78684 162176 78736
rect 164516 78684 164568 78736
rect 166540 78684 166592 78736
rect 168656 78684 168708 78736
rect 554780 78684 554832 78736
rect 157892 78616 157944 78668
rect 158076 78616 158128 78668
rect 160560 78616 160612 78668
rect 160836 78616 160888 78668
rect 160928 78616 160980 78668
rect 170864 78616 170916 78668
rect 139676 78548 139728 78600
rect 171784 78616 171836 78668
rect 171968 78616 172020 78668
rect 179420 78616 179472 78668
rect 172428 78548 172480 78600
rect 173624 78548 173676 78600
rect 128636 78480 128688 78532
rect 131212 78480 131264 78532
rect 140780 78480 140832 78532
rect 166908 78480 166960 78532
rect 142620 78412 142672 78464
rect 160928 78412 160980 78464
rect 161204 78412 161256 78464
rect 163136 78412 163188 78464
rect 171692 78480 171744 78532
rect 172060 78480 172112 78532
rect 178960 78548 179012 78600
rect 125324 78344 125376 78396
rect 125600 78344 125652 78396
rect 142252 78344 142304 78396
rect 171232 78412 171284 78464
rect 175188 78412 175240 78464
rect 164792 78344 164844 78396
rect 167000 78344 167052 78396
rect 167092 78344 167144 78396
rect 173164 78344 173216 78396
rect 120816 78276 120868 78328
rect 129096 78276 129148 78328
rect 131212 78276 131264 78328
rect 131948 78276 132000 78328
rect 152648 78276 152700 78328
rect 160928 78276 160980 78328
rect 161112 78276 161164 78328
rect 247684 78276 247736 78328
rect 125232 78208 125284 78260
rect 132960 78208 133012 78260
rect 154212 78208 154264 78260
rect 154672 78208 154724 78260
rect 160744 78208 160796 78260
rect 161296 78208 161348 78260
rect 162400 78208 162452 78260
rect 253204 78208 253256 78260
rect 89720 78140 89772 78192
rect 132408 78140 132460 78192
rect 133972 78140 134024 78192
rect 134432 78140 134484 78192
rect 155132 78140 155184 78192
rect 161020 78140 161072 78192
rect 162952 78140 163004 78192
rect 163596 78140 163648 78192
rect 165344 78140 165396 78192
rect 168748 78140 168800 78192
rect 170128 78140 170180 78192
rect 170680 78140 170732 78192
rect 171048 78140 171100 78192
rect 322204 78140 322256 78192
rect 57244 78072 57296 78124
rect 126980 78072 127032 78124
rect 140872 78072 140924 78124
rect 159640 78072 159692 78124
rect 162124 78072 162176 78124
rect 162308 78072 162360 78124
rect 471980 78072 472032 78124
rect 46204 78004 46256 78056
rect 126336 78004 126388 78056
rect 129096 78004 129148 78056
rect 129464 78004 129516 78056
rect 129648 78004 129700 78056
rect 129832 78004 129884 78056
rect 134432 78004 134484 78056
rect 135168 78004 135220 78056
rect 140320 78004 140372 78056
rect 148692 78004 148744 78056
rect 150256 78004 150308 78056
rect 154304 78004 154356 78056
rect 162400 78004 162452 78056
rect 162768 78004 162820 78056
rect 480260 78004 480312 78056
rect 22744 77936 22796 77988
rect 122932 77936 122984 77988
rect 125140 77936 125192 77988
rect 127072 77936 127124 77988
rect 129004 77936 129056 77988
rect 131396 77936 131448 77988
rect 132224 77936 132276 77988
rect 132684 77936 132736 77988
rect 133880 77936 133932 77988
rect 135904 77936 135956 77988
rect 156144 77936 156196 77988
rect 125324 77868 125376 77920
rect 133420 77868 133472 77920
rect 135444 77868 135496 77920
rect 136548 77868 136600 77920
rect 160652 77936 160704 77988
rect 162308 77868 162360 77920
rect 163228 77868 163280 77920
rect 164056 77868 164108 77920
rect 164792 77868 164844 77920
rect 165160 77868 165212 77920
rect 168748 77936 168800 77988
rect 498200 77936 498252 77988
rect 180064 77868 180116 77920
rect 126980 77800 127032 77852
rect 129372 77800 129424 77852
rect 129740 77800 129792 77852
rect 130568 77800 130620 77852
rect 133052 77800 133104 77852
rect 133236 77800 133288 77852
rect 151544 77800 151596 77852
rect 156144 77800 156196 77852
rect 158628 77800 158680 77852
rect 174544 77800 174596 77852
rect 123484 77732 123536 77784
rect 134892 77732 134944 77784
rect 159272 77732 159324 77784
rect 175924 77732 175976 77784
rect 122564 77664 122616 77716
rect 127624 77664 127676 77716
rect 132776 77664 132828 77716
rect 133236 77664 133288 77716
rect 138020 77664 138072 77716
rect 139032 77664 139084 77716
rect 139308 77664 139360 77716
rect 129372 77596 129424 77648
rect 130200 77596 130252 77648
rect 143632 77596 143684 77648
rect 153292 77596 153344 77648
rect 131672 77528 131724 77580
rect 132040 77528 132092 77580
rect 136640 77528 136692 77580
rect 139032 77528 139084 77580
rect 130016 77460 130068 77512
rect 135628 77460 135680 77512
rect 147772 77460 147824 77512
rect 158352 77664 158404 77716
rect 172428 77664 172480 77716
rect 159916 77596 159968 77648
rect 171416 77596 171468 77648
rect 160376 77528 160428 77580
rect 160652 77528 160704 77580
rect 171600 77528 171652 77580
rect 580632 77528 580684 77580
rect 126336 77392 126388 77444
rect 130384 77392 130436 77444
rect 133512 77392 133564 77444
rect 136916 77392 136968 77444
rect 149704 77392 149756 77444
rect 152648 77392 152700 77444
rect 167460 77460 167512 77512
rect 168288 77460 168340 77512
rect 171784 77460 171836 77512
rect 158260 77392 158312 77444
rect 171324 77392 171376 77444
rect 171692 77392 171744 77444
rect 144920 77324 144972 77376
rect 162216 77324 162268 77376
rect 163412 77324 163464 77376
rect 172060 77324 172112 77376
rect 142436 77256 142488 77308
rect 142804 77256 142856 77308
rect 148876 77256 148928 77308
rect 148968 77188 149020 77240
rect 149520 77188 149572 77240
rect 151268 77256 151320 77308
rect 156144 77256 156196 77308
rect 157064 77256 157116 77308
rect 153016 77188 153068 77240
rect 154212 77188 154264 77240
rect 178776 77188 178828 77240
rect 527180 77188 527232 77240
rect 120908 77120 120960 77172
rect 171876 77120 171928 77172
rect 121000 77052 121052 77104
rect 172612 77052 172664 77104
rect 153844 76984 153896 77036
rect 211804 76984 211856 77036
rect 152372 76916 152424 76968
rect 226340 76916 226392 76968
rect 124864 76848 124916 76900
rect 134800 76848 134852 76900
rect 146944 76848 146996 76900
rect 240140 76848 240192 76900
rect 102140 76780 102192 76832
rect 132500 76780 132552 76832
rect 135628 76780 135680 76832
rect 135812 76780 135864 76832
rect 145656 76780 145708 76832
rect 260840 76780 260892 76832
rect 86960 76712 87012 76764
rect 132316 76712 132368 76764
rect 148324 76712 148376 76764
rect 69020 76644 69072 76696
rect 128544 76644 128596 76696
rect 132592 76644 132644 76696
rect 133144 76644 133196 76696
rect 145472 76644 145524 76696
rect 145656 76644 145708 76696
rect 150532 76644 150584 76696
rect 153016 76712 153068 76764
rect 288440 76712 288492 76764
rect 44180 76576 44232 76628
rect 128360 76576 128412 76628
rect 143172 76576 143224 76628
rect 152372 76576 152424 76628
rect 296720 76644 296772 76696
rect 324412 76576 324464 76628
rect 30380 76508 30432 76560
rect 127900 76508 127952 76560
rect 137376 76508 137428 76560
rect 144552 76508 144604 76560
rect 152096 76508 152148 76560
rect 152280 76508 152332 76560
rect 158720 76508 158772 76560
rect 159272 76508 159324 76560
rect 159456 76508 159508 76560
rect 160008 76508 160060 76560
rect 160192 76508 160244 76560
rect 454040 76508 454092 76560
rect 122840 76440 122892 76492
rect 135076 76440 135128 76492
rect 150256 76440 150308 76492
rect 197360 76440 197412 76492
rect 119988 76372 120040 76424
rect 172888 76372 172940 76424
rect 127624 76304 127676 76356
rect 129188 76304 129240 76356
rect 156052 76304 156104 76356
rect 156420 76304 156472 76356
rect 158720 76304 158772 76356
rect 159732 76304 159784 76356
rect 127256 76236 127308 76288
rect 128268 76236 128320 76288
rect 151820 76236 151872 76288
rect 152280 76236 152332 76288
rect 155776 76236 155828 76288
rect 159640 76236 159692 76288
rect 143632 76168 143684 76220
rect 144092 76168 144144 76220
rect 154580 76168 154632 76220
rect 155132 76168 155184 76220
rect 154672 76100 154724 76152
rect 155224 76100 155276 76152
rect 143816 76032 143868 76084
rect 143908 76032 143960 76084
rect 144092 76032 144144 76084
rect 153476 76032 153528 76084
rect 155868 76032 155920 76084
rect 156236 76032 156288 76084
rect 156512 76032 156564 76084
rect 125508 75896 125560 75948
rect 126244 75896 126296 75948
rect 127440 75896 127492 75948
rect 127716 75896 127768 75948
rect 141056 75896 141108 75948
rect 141700 75896 141752 75948
rect 142160 75896 142212 75948
rect 143080 75896 143132 75948
rect 143908 75896 143960 75948
rect 153384 75896 153436 75948
rect 154120 75896 154172 75948
rect 154580 75896 154632 75948
rect 155500 75896 155552 75948
rect 157248 75896 157300 75948
rect 158260 75896 158312 75948
rect 122104 75828 122156 75880
rect 127348 75828 127400 75880
rect 153292 75828 153344 75880
rect 153568 75828 153620 75880
rect 155960 75828 156012 75880
rect 156604 75828 156656 75880
rect 120724 75760 120776 75812
rect 128452 75760 128504 75812
rect 154764 75760 154816 75812
rect 155040 75760 155092 75812
rect 156788 75760 156840 75812
rect 127348 75692 127400 75744
rect 128176 75692 128228 75744
rect 129832 75692 129884 75744
rect 130016 75692 130068 75744
rect 142252 75692 142304 75744
rect 142988 75692 143040 75744
rect 151820 75692 151872 75744
rect 152188 75692 152240 75744
rect 122288 75624 122340 75676
rect 128084 75624 128136 75676
rect 158996 75624 159048 75676
rect 130016 75556 130068 75608
rect 130660 75556 130712 75608
rect 159916 75556 159968 75608
rect 166724 75556 166776 75608
rect 122196 75488 122248 75540
rect 130476 75488 130528 75540
rect 154764 75488 154816 75540
rect 155408 75488 155460 75540
rect 162216 75488 162268 75540
rect 396080 75556 396132 75608
rect 121460 75420 121512 75472
rect 134984 75420 135036 75472
rect 136824 75420 136876 75472
rect 137652 75420 137704 75472
rect 163964 75420 164016 75472
rect 51080 75352 51132 75404
rect 129096 75352 129148 75404
rect 136916 75352 136968 75404
rect 137284 75352 137336 75404
rect 149336 75352 149388 75404
rect 149520 75352 149572 75404
rect 155960 75352 156012 75404
rect 156696 75352 156748 75404
rect 164424 75352 164476 75404
rect 164700 75352 164752 75404
rect 165804 75352 165856 75404
rect 166540 75352 166592 75404
rect 107660 75284 107712 75336
rect 131580 75284 131632 75336
rect 132684 75284 132736 75336
rect 133604 75284 133656 75336
rect 135444 75284 135496 75336
rect 136180 75284 136232 75336
rect 144920 75284 144972 75336
rect 145840 75284 145892 75336
rect 146208 75284 146260 75336
rect 146852 75284 146904 75336
rect 147680 75284 147732 75336
rect 148600 75284 148652 75336
rect 151912 75284 151964 75336
rect 152372 75284 152424 75336
rect 164608 75284 164660 75336
rect 431960 75488 432012 75540
rect 166816 75420 166868 75472
rect 438860 75420 438912 75472
rect 467840 75352 467892 75404
rect 42800 75216 42852 75268
rect 128360 75216 128412 75268
rect 128728 75216 128780 75268
rect 129648 75216 129700 75268
rect 130292 75216 130344 75268
rect 131028 75216 131080 75268
rect 132868 75216 132920 75268
rect 133696 75216 133748 75268
rect 134248 75216 134300 75268
rect 134708 75216 134760 75268
rect 135904 75216 135956 75268
rect 136364 75216 136416 75268
rect 136824 75216 136876 75268
rect 137468 75216 137520 75268
rect 138112 75216 138164 75268
rect 138664 75216 138716 75268
rect 139676 75216 139728 75268
rect 140136 75216 140188 75268
rect 144000 75216 144052 75268
rect 144460 75216 144512 75268
rect 145380 75216 145432 75268
rect 145748 75216 145800 75268
rect 146484 75216 146536 75268
rect 146760 75216 146812 75268
rect 146944 75216 146996 75268
rect 147128 75216 147180 75268
rect 148048 75216 148100 75268
rect 148416 75216 148468 75268
rect 149336 75216 149388 75268
rect 149888 75216 149940 75268
rect 150716 75216 150768 75268
rect 151084 75216 151136 75268
rect 152188 75216 152240 75268
rect 152556 75216 152608 75268
rect 153200 75216 153252 75268
rect 153936 75216 153988 75268
rect 157524 75216 157576 75268
rect 158076 75216 158128 75268
rect 160376 75216 160428 75268
rect 160744 75216 160796 75268
rect 161572 75216 161624 75268
rect 162032 75216 162084 75268
rect 163044 75216 163096 75268
rect 163412 75216 163464 75268
rect 164700 75216 164752 75268
rect 164976 75216 165028 75268
rect 165804 75216 165856 75268
rect 166356 75216 166408 75268
rect 490012 75284 490064 75336
rect 499580 75216 499632 75268
rect 6920 75148 6972 75200
rect 123024 75148 123076 75200
rect 128544 75148 128596 75200
rect 128912 75148 128964 75200
rect 132960 75148 133012 75200
rect 133788 75148 133840 75200
rect 135536 75148 135588 75200
rect 136272 75148 136324 75200
rect 137008 75148 137060 75200
rect 137192 75148 137244 75200
rect 139952 75148 140004 75200
rect 140228 75148 140280 75200
rect 145104 75148 145156 75200
rect 145472 75148 145524 75200
rect 146576 75148 146628 75200
rect 146852 75148 146904 75200
rect 147772 75148 147824 75200
rect 148508 75148 148560 75200
rect 151912 75148 151964 75200
rect 152924 75148 152976 75200
rect 157800 75148 157852 75200
rect 158168 75148 158220 75200
rect 160192 75148 160244 75200
rect 160836 75148 160888 75200
rect 162860 75148 162912 75200
rect 163504 75148 163556 75200
rect 164608 75148 164660 75200
rect 165160 75148 165212 75200
rect 167460 75148 167512 75200
rect 167828 75148 167880 75200
rect 168380 75148 168432 75200
rect 168748 75148 168800 75200
rect 168840 75148 168892 75200
rect 169392 75148 169444 75200
rect 169760 75148 169812 75200
rect 170312 75148 170364 75200
rect 173992 75148 174044 75200
rect 174360 75148 174412 75200
rect 128636 75080 128688 75132
rect 129280 75080 129332 75132
rect 135720 75080 135772 75132
rect 136456 75080 136508 75132
rect 138756 75080 138808 75132
rect 140412 75080 140464 75132
rect 141240 75080 141292 75132
rect 141516 75080 141568 75132
rect 142528 75080 142580 75132
rect 142804 75080 142856 75132
rect 146484 75080 146536 75132
rect 147496 75080 147548 75132
rect 150716 75080 150768 75132
rect 151360 75080 151412 75132
rect 161572 75080 161624 75132
rect 162124 75080 162176 75132
rect 163044 75080 163096 75132
rect 163872 75080 163924 75132
rect 167092 75080 167144 75132
rect 167920 75080 167972 75132
rect 170220 75080 170272 75132
rect 170864 75080 170916 75132
rect 128360 75012 128412 75064
rect 136548 75012 136600 75064
rect 137008 75012 137060 75064
rect 137744 75012 137796 75064
rect 145104 75012 145156 75064
rect 145932 75012 145984 75064
rect 146576 75012 146628 75064
rect 147220 75012 147272 75064
rect 168380 75012 168432 75064
rect 168564 75012 168616 75064
rect 169760 75012 169812 75064
rect 170496 75012 170548 75064
rect 140964 74944 141016 74996
rect 141792 74944 141844 74996
rect 169576 74944 169628 74996
rect 564440 75148 564492 75200
rect 131672 74876 131724 74928
rect 132132 74876 132184 74928
rect 146300 74876 146352 74928
rect 147220 74876 147272 74928
rect 168564 74876 168616 74928
rect 169116 74876 169168 74928
rect 124772 74808 124824 74860
rect 125416 74808 125468 74860
rect 167000 74468 167052 74520
rect 173348 74468 173400 74520
rect 141976 74196 142028 74248
rect 209780 74196 209832 74248
rect 144828 74128 144880 74180
rect 216680 74128 216732 74180
rect 118700 74060 118752 74112
rect 134064 74060 134116 74112
rect 143448 74060 143500 74112
rect 223580 74060 223632 74112
rect 93952 73992 94004 74044
rect 133236 73992 133288 74044
rect 145656 73992 145708 74044
rect 251180 73992 251232 74044
rect 64880 73924 64932 73976
rect 129740 73924 129792 73976
rect 152648 73924 152700 73976
rect 318800 73924 318852 73976
rect 27620 73856 27672 73908
rect 126888 73856 126940 73908
rect 153108 73856 153160 73908
rect 354680 73856 354732 73908
rect 26240 73788 26292 73840
rect 122564 73788 122616 73840
rect 161020 73788 161072 73840
rect 375380 73788 375432 73840
rect 137560 73176 137612 73228
rect 142988 73176 143040 73228
rect 170956 73108 171008 73160
rect 580172 73108 580224 73160
rect 126428 72768 126480 72820
rect 126796 72768 126848 72820
rect 140872 72700 140924 72752
rect 141424 72700 141476 72752
rect 148968 72632 149020 72684
rect 291200 72632 291252 72684
rect 149060 72564 149112 72616
rect 311900 72564 311952 72616
rect 152740 72496 152792 72548
rect 340880 72496 340932 72548
rect 155868 72428 155920 72480
rect 357440 72428 357492 72480
rect 165068 72360 165120 72412
rect 171876 72360 171928 72412
rect 3424 71680 3476 71732
rect 179604 71680 179656 71732
rect 78680 71000 78732 71052
rect 132040 71000 132092 71052
rect 138940 71000 138992 71052
rect 152556 71000 152608 71052
rect 158352 71000 158404 71052
rect 284392 71000 284444 71052
rect 138664 70320 138716 70372
rect 142804 70320 142856 70372
rect 141516 70048 141568 70100
rect 209872 70048 209924 70100
rect 155316 69980 155368 70032
rect 382280 69980 382332 70032
rect 156604 69912 156656 69964
rect 390560 69912 390612 69964
rect 171692 69844 171744 69896
rect 426440 69844 426492 69896
rect 164884 69776 164936 69828
rect 505100 69776 505152 69828
rect 166540 69708 166592 69760
rect 518900 69708 518952 69760
rect 170312 69640 170364 69692
rect 568580 69640 568632 69692
rect 170220 68960 170272 69012
rect 171692 68960 171744 69012
rect 140044 68620 140096 68672
rect 184940 68620 184992 68672
rect 142712 68552 142764 68604
rect 218060 68552 218112 68604
rect 157064 68484 157116 68536
rect 320180 68484 320232 68536
rect 153752 68416 153804 68468
rect 362960 68416 363012 68468
rect 159272 68348 159324 68400
rect 427820 68348 427872 68400
rect 169484 68280 169536 68332
rect 564532 68280 564584 68332
rect 139952 67396 140004 67448
rect 189080 67396 189132 67448
rect 147220 67328 147272 67380
rect 270500 67328 270552 67380
rect 149704 67260 149756 67312
rect 306380 67260 306432 67312
rect 160836 67192 160888 67244
rect 347780 67192 347832 67244
rect 152464 67124 152516 67176
rect 340972 67124 341024 67176
rect 159180 67056 159232 67108
rect 437480 67056 437532 67108
rect 162032 66988 162084 67040
rect 462320 66988 462372 67040
rect 167736 66920 167788 66972
rect 539600 66920 539652 66972
rect 167644 66852 167696 66904
rect 543740 66852 543792 66904
rect 137284 66172 137336 66224
rect 140044 66172 140096 66224
rect 138572 66104 138624 66156
rect 141516 66104 141568 66156
rect 141332 65900 141384 65952
rect 202880 65900 202932 65952
rect 141424 65832 141476 65884
rect 207020 65832 207072 65884
rect 142620 65764 142672 65816
rect 220820 65764 220872 65816
rect 145472 65696 145524 65748
rect 251272 65696 251324 65748
rect 145564 65628 145616 65680
rect 256700 65628 256752 65680
rect 153660 65560 153712 65612
rect 358820 65560 358872 65612
rect 102232 65492 102284 65544
rect 125324 65492 125376 65544
rect 155224 65492 155276 65544
rect 376760 65492 376812 65544
rect 144276 64472 144328 64524
rect 234620 64472 234672 64524
rect 144184 64404 144236 64456
rect 238760 64404 238812 64456
rect 148232 64336 148284 64388
rect 292580 64336 292632 64388
rect 152372 64268 152424 64320
rect 338120 64268 338172 64320
rect 162584 64200 162636 64252
rect 368480 64200 368532 64252
rect 169024 64132 169076 64184
rect 561680 64132 561732 64184
rect 147036 63112 147088 63164
rect 274640 63112 274692 63164
rect 149612 63044 149664 63096
rect 309140 63044 309192 63096
rect 155132 62976 155184 63028
rect 374000 62976 374052 63028
rect 157984 62908 158036 62960
rect 408500 62908 408552 62960
rect 163596 62840 163648 62892
rect 488540 62840 488592 62892
rect 168932 62772 168984 62824
rect 557540 62772 557592 62824
rect 139860 61480 139912 61532
rect 185032 61480 185084 61532
rect 157892 61412 157944 61464
rect 412640 61412 412692 61464
rect 166356 61344 166408 61396
rect 525800 61344 525852 61396
rect 118516 60664 118568 60716
rect 580172 60664 580224 60716
rect 137192 59984 137244 60036
rect 138664 59984 138716 60036
rect 159088 59984 159140 60036
rect 433340 59984 433392 60036
rect 156512 58624 156564 58676
rect 401600 58624 401652 58676
rect 163504 57264 163556 57316
rect 481640 57264 481692 57316
rect 164792 57196 164844 57248
rect 507860 57196 507912 57248
rect 95240 53048 95292 53100
rect 125232 53048 125284 53100
rect 182824 46860 182876 46912
rect 580172 46860 580224 46912
rect 139768 46180 139820 46232
rect 180800 46180 180852 46232
rect 3424 45500 3476 45552
rect 174084 45500 174136 45552
rect 135996 44956 136048 45008
rect 142620 44956 142672 45008
rect 70400 44888 70452 44940
rect 130292 44888 130344 44940
rect 34520 44820 34572 44872
rect 127348 44820 127400 44872
rect 138480 44820 138532 44872
rect 147036 44820 147088 44872
rect 171600 43392 171652 43444
rect 411260 43392 411312 43444
rect 19340 42032 19392 42084
rect 125140 42032 125192 42084
rect 162216 42032 162268 42084
rect 390652 42032 390704 42084
rect 172428 40672 172480 40724
rect 418160 40672 418212 40724
rect 120080 40264 120132 40316
rect 123484 40264 123536 40316
rect 172336 39312 172388 39364
rect 404360 39312 404412 39364
rect 172244 37884 172296 37936
rect 397460 37884 397512 37936
rect 88340 36524 88392 36576
rect 125048 36524 125100 36576
rect 145380 35572 145432 35624
rect 259460 35572 259512 35624
rect 146944 35504 146996 35556
rect 276020 35504 276072 35556
rect 148140 35436 148192 35488
rect 287060 35436 287112 35488
rect 148048 35368 148100 35420
rect 293960 35368 294012 35420
rect 149520 35300 149572 35352
rect 305000 35300 305052 35352
rect 149428 35232 149480 35284
rect 307760 35232 307812 35284
rect 159732 35164 159784 35216
rect 382372 35164 382424 35216
rect 139676 34076 139728 34128
rect 187700 34076 187752 34128
rect 141148 34008 141200 34060
rect 198740 34008 198792 34060
rect 141056 33940 141108 33992
rect 201500 33940 201552 33992
rect 141240 33872 141292 33924
rect 205640 33872 205692 33924
rect 144092 33804 144144 33856
rect 234712 33804 234764 33856
rect 146852 33736 146904 33788
rect 269120 33736 269172 33788
rect 171692 33056 171744 33108
rect 580172 33056 580224 33108
rect 3424 32988 3476 33040
rect 180892 32988 180944 33040
rect 156420 32716 156472 32768
rect 391940 32716 391992 32768
rect 160008 32648 160060 32700
rect 434720 32648 434772 32700
rect 161940 32580 161992 32632
rect 463700 32580 463752 32632
rect 163412 32512 163464 32564
rect 481732 32512 481784 32564
rect 167552 32444 167604 32496
rect 539692 32444 539744 32496
rect 170128 32376 170180 32428
rect 574100 32376 574152 32428
rect 144000 31424 144052 31476
rect 242900 31424 242952 31476
rect 146760 31356 146812 31408
rect 267832 31356 267884 31408
rect 147956 31288 148008 31340
rect 289820 31288 289872 31340
rect 154120 31220 154172 31272
rect 332600 31220 332652 31272
rect 153568 31152 153620 31204
rect 357532 31152 357584 31204
rect 156972 31084 157024 31136
rect 389180 31084 389232 31136
rect 166264 31016 166316 31068
rect 524420 31016 524472 31068
rect 140872 30064 140924 30116
rect 204260 30064 204312 30116
rect 140964 29996 141016 30048
rect 208400 29996 208452 30048
rect 143908 29928 143960 29980
rect 233240 29928 233292 29980
rect 143816 29860 143868 29912
rect 236000 29860 236052 29912
rect 145288 29792 145340 29844
rect 253940 29792 253992 29844
rect 145196 29724 145248 29776
rect 258080 29724 258132 29776
rect 166172 29656 166224 29708
rect 521660 29656 521712 29708
rect 167460 29588 167512 29640
rect 542360 29588 542412 29640
rect 148692 28500 148744 28552
rect 190460 28500 190512 28552
rect 139584 28432 139636 28484
rect 186320 28432 186372 28484
rect 140780 28364 140832 28416
rect 201592 28364 201644 28416
rect 146668 28296 146720 28348
rect 271880 28296 271932 28348
rect 147864 28228 147916 28280
rect 285680 28228 285732 28280
rect 322204 28228 322256 28280
rect 581000 28228 581052 28280
rect 140504 27276 140556 27328
rect 176752 27276 176804 27328
rect 139400 27208 139452 27260
rect 179420 27208 179472 27260
rect 139492 27140 139544 27192
rect 183560 27140 183612 27192
rect 146576 27072 146628 27124
rect 276112 27072 276164 27124
rect 149336 27004 149388 27056
rect 310520 27004 310572 27056
rect 152280 26936 152332 26988
rect 339500 26936 339552 26988
rect 164700 26868 164752 26920
rect 506480 26868 506532 26920
rect 142528 25984 142580 26036
rect 222200 25984 222252 26036
rect 146484 25916 146536 25968
rect 278780 25916 278832 25968
rect 149244 25848 149296 25900
rect 307852 25848 307904 25900
rect 152188 25780 152240 25832
rect 346400 25780 346452 25832
rect 166080 25712 166132 25764
rect 517520 25712 517572 25764
rect 170680 25644 170732 25696
rect 558920 25644 558972 25696
rect 168840 25576 168892 25628
rect 563060 25576 563112 25628
rect 170036 25508 170088 25560
rect 572720 25508 572772 25560
rect 142344 24556 142396 24608
rect 215300 24556 215352 24608
rect 142436 24488 142488 24540
rect 218152 24488 218204 24540
rect 147772 24420 147824 24472
rect 292672 24420 292724 24472
rect 155040 24352 155092 24404
rect 374092 24352 374144 24404
rect 167368 24284 167420 24336
rect 467104 24284 467156 24336
rect 167276 24216 167328 24268
rect 535460 24216 535512 24268
rect 167184 24148 167236 24200
rect 538220 24148 538272 24200
rect 168748 24080 168800 24132
rect 552020 24080 552072 24132
rect 149152 23332 149204 23384
rect 303620 23332 303672 23384
rect 3424 23264 3476 23316
rect 173992 23264 174044 23316
rect 153476 23196 153528 23248
rect 360200 23196 360252 23248
rect 154948 23128 155000 23180
rect 379520 23128 379572 23180
rect 164516 23060 164568 23112
rect 498292 23060 498344 23112
rect 164608 22992 164660 23044
rect 509240 22992 509292 23044
rect 165896 22924 165948 22976
rect 516140 22924 516192 22976
rect 165988 22856 166040 22908
rect 520280 22856 520332 22908
rect 74540 22788 74592 22840
rect 128452 22788 128504 22840
rect 168656 22788 168708 22840
rect 556160 22788 556212 22840
rect 118424 22720 118476 22772
rect 580172 22720 580224 22772
rect 152096 21632 152148 21684
rect 343640 21632 343692 21684
rect 160652 21564 160704 21616
rect 447140 21564 447192 21616
rect 161848 21496 161900 21548
rect 473360 21496 473412 21548
rect 163320 21428 163372 21480
rect 484400 21428 484452 21480
rect 124312 21360 124364 21412
rect 134340 21360 134392 21412
rect 164424 21360 164476 21412
rect 506572 21360 506624 21412
rect 145012 20340 145064 20392
rect 255320 20340 255372 20392
rect 145104 20272 145156 20324
rect 262220 20272 262272 20324
rect 146392 20204 146444 20256
rect 273260 20204 273312 20256
rect 247684 20136 247736 20188
rect 456800 20136 456852 20188
rect 138388 20068 138440 20120
rect 162860 20068 162912 20120
rect 253204 20068 253256 20120
rect 465080 20068 465132 20120
rect 85580 20000 85632 20052
rect 131672 20000 131724 20052
rect 160560 20000 160612 20052
rect 455420 20000 455472 20052
rect 45560 19932 45612 19984
rect 120816 19932 120868 19984
rect 161756 19932 161808 19984
rect 465172 19932 465224 19984
rect 160468 18844 160520 18896
rect 448520 18844 448572 18896
rect 160376 18776 160428 18828
rect 451280 18776 451332 18828
rect 117320 18708 117372 18760
rect 134248 18708 134300 18760
rect 168472 18708 168524 18760
rect 553400 18708 553452 18760
rect 31760 18640 31812 18692
rect 122288 18640 122340 18692
rect 168380 18640 168432 18692
rect 556252 18640 556304 18692
rect 4160 18572 4212 18624
rect 126244 18572 126296 18624
rect 168564 18572 168616 18624
rect 560300 18572 560352 18624
rect 157708 17552 157760 17604
rect 415400 17552 415452 17604
rect 157800 17484 157852 17536
rect 419540 17484 419592 17536
rect 171968 17416 172020 17468
rect 440240 17416 440292 17468
rect 160284 17348 160336 17400
rect 448612 17348 448664 17400
rect 163228 17280 163280 17332
rect 492680 17280 492732 17332
rect 167092 17212 167144 17264
rect 545120 17212 545172 17264
rect 154856 16124 154908 16176
rect 378416 16124 378468 16176
rect 156328 16056 156380 16108
rect 395344 16056 395396 16108
rect 156236 15988 156288 16040
rect 398840 15988 398892 16040
rect 174544 15920 174596 15972
rect 425704 15920 425756 15972
rect 14280 15852 14332 15904
rect 124956 15852 125008 15904
rect 167920 15852 167972 15904
rect 541992 15852 542044 15904
rect 143724 14764 143776 14816
rect 241704 14764 241756 14816
rect 154672 14696 154724 14748
rect 381176 14696 381228 14748
rect 154764 14628 154816 14680
rect 384304 14628 384356 14680
rect 154580 14560 154632 14612
rect 385960 14560 386012 14612
rect 114008 14492 114060 14544
rect 134156 14492 134208 14544
rect 158904 14492 158956 14544
rect 436744 14492 436796 14544
rect 39120 14424 39172 14476
rect 120724 14424 120776 14476
rect 164332 14424 164384 14476
rect 502984 14424 503036 14476
rect 152004 13404 152056 13456
rect 345296 13404 345348 13456
rect 151912 13336 151964 13388
rect 349160 13336 349212 13388
rect 153384 13268 153436 13320
rect 365720 13268 365772 13320
rect 157616 13200 157668 13252
rect 417424 13200 417476 13252
rect 158812 13132 158864 13184
rect 429200 13132 429252 13184
rect 160192 13064 160244 13116
rect 453304 13064 453356 13116
rect 143632 11976 143684 12028
rect 237656 11976 237708 12028
rect 150348 11908 150400 11960
rect 313832 11908 313884 11960
rect 135812 11840 135864 11892
rect 157432 11840 157484 11892
rect 414296 11840 414348 11892
rect 135720 11636 135772 11688
rect 157524 11772 157576 11824
rect 415492 11772 415544 11824
rect 165804 11704 165856 11756
rect 523776 11704 523828 11756
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 184940 11636 184992 11688
rect 186136 11636 186188 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 106464 10616 106516 10668
rect 132960 10616 133012 10668
rect 99840 10548 99892 10600
rect 133052 10548 133104 10600
rect 147680 10548 147732 10600
rect 295616 10548 295668 10600
rect 81624 10480 81676 10532
rect 131580 10480 131632 10532
rect 154488 10480 154540 10532
rect 364616 10480 364668 10532
rect 35992 10412 36044 10464
rect 127256 10412 127308 10464
rect 156052 10412 156104 10464
rect 394240 10412 394292 10464
rect 28448 10344 28500 10396
rect 127164 10344 127216 10396
rect 156144 10344 156196 10396
rect 398932 10344 398984 10396
rect 11152 10276 11204 10328
rect 126152 10276 126204 10328
rect 163136 10276 163188 10328
rect 486424 10276 486476 10328
rect 67916 9324 67968 9376
rect 130200 9324 130252 9376
rect 64328 9256 64380 9308
rect 126336 9256 126388 9308
rect 144920 9256 144972 9308
rect 260656 9256 260708 9308
rect 63224 9188 63276 9240
rect 130108 9188 130160 9240
rect 146300 9188 146352 9240
rect 278320 9188 278372 9240
rect 60832 9120 60884 9172
rect 129096 9120 129148 9172
rect 151820 9120 151872 9172
rect 343364 9120 343416 9172
rect 53748 9052 53800 9104
rect 128728 9052 128780 9104
rect 161664 9052 161716 9104
rect 471060 9052 471112 9104
rect 50160 8984 50212 9036
rect 126980 8984 127032 9036
rect 163044 8984 163096 9036
rect 492312 8984 492364 9036
rect 572 8916 624 8968
rect 124220 8916 124272 8968
rect 169944 8916 169996 8968
rect 571524 8916 571576 8968
rect 116400 7896 116452 7948
rect 134064 7896 134116 7948
rect 142252 7896 142304 7948
rect 225144 7896 225196 7948
rect 105728 7828 105780 7880
rect 132868 7828 132920 7880
rect 143540 7828 143592 7880
rect 242992 7828 243044 7880
rect 98644 7760 98696 7812
rect 132776 7760 132828 7812
rect 155960 7760 156012 7812
rect 401324 7760 401376 7812
rect 48964 7692 49016 7744
rect 128636 7692 128688 7744
rect 160100 7692 160152 7744
rect 446220 7692 446272 7744
rect 44272 7624 44324 7676
rect 128544 7624 128596 7676
rect 161572 7624 161624 7676
rect 469864 7624 469916 7676
rect 9956 7556 10008 7608
rect 126060 7556 126112 7608
rect 164240 7556 164292 7608
rect 504180 7556 504232 7608
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 151084 6740 151136 6792
rect 323308 6740 323360 6792
rect 150900 6672 150952 6724
rect 326804 6672 326856 6724
rect 115204 6604 115256 6656
rect 134708 6604 134760 6656
rect 150992 6604 151044 6656
rect 329196 6604 329248 6656
rect 104532 6536 104584 6588
rect 132684 6536 132736 6588
rect 150808 6536 150860 6588
rect 330392 6536 330444 6588
rect 84476 6468 84528 6520
rect 131304 6468 131356 6520
rect 157340 6468 157392 6520
rect 410800 6468 410852 6520
rect 80888 6400 80940 6452
rect 131488 6400 131540 6452
rect 175924 6400 175976 6452
rect 433248 6400 433300 6452
rect 77392 6332 77444 6384
rect 131396 6332 131448 6384
rect 158720 6332 158772 6384
rect 441528 6332 441580 6384
rect 25320 6264 25372 6316
rect 57244 6264 57296 6316
rect 66720 6264 66772 6316
rect 130016 6264 130068 6316
rect 161480 6264 161532 6316
rect 467472 6264 467524 6316
rect 33600 6196 33652 6248
rect 127532 6196 127584 6248
rect 140412 6196 140464 6248
rect 156604 6196 156656 6248
rect 169852 6196 169904 6248
rect 572720 6196 572772 6248
rect 18236 6128 18288 6180
rect 125968 6128 126020 6180
rect 138296 6128 138348 6180
rect 162492 6128 162544 6180
rect 169760 6128 169812 6180
rect 576308 6128 576360 6180
rect 101036 5312 101088 5364
rect 133144 5312 133196 5364
rect 97448 5244 97500 5296
rect 132592 5244 132644 5296
rect 86868 5176 86920 5228
rect 132040 5176 132092 5228
rect 138112 5176 138164 5228
rect 169576 5176 169628 5228
rect 15936 5040 15988 5092
rect 59636 5108 59688 5160
rect 129924 5108 129976 5160
rect 142160 5108 142212 5160
rect 220452 5108 220504 5160
rect 46204 5040 46256 5092
rect 52552 5040 52604 5092
rect 129648 5040 129700 5092
rect 137100 5040 137152 5092
rect 148324 5040 148376 5092
rect 153292 5040 153344 5092
rect 365812 5040 365864 5092
rect 33232 4972 33284 5024
rect 127440 4972 127492 5024
rect 138020 4972 138072 5024
rect 171968 4972 172020 5024
rect 180064 4972 180116 5024
rect 450912 4972 450964 5024
rect 6460 4904 6512 4956
rect 22744 4904 22796 4956
rect 24216 4904 24268 4956
rect 122104 4904 122156 4956
rect 136916 4904 136968 4956
rect 150624 4904 150676 4956
rect 162952 4904 163004 4956
rect 487620 4904 487672 4956
rect 13544 4836 13596 4888
rect 125876 4836 125928 4888
rect 137008 4836 137060 4888
rect 157800 4836 157852 4888
rect 165620 4836 165672 4888
rect 523040 4836 523092 4888
rect 8760 4768 8812 4820
rect 125784 4768 125836 4820
rect 138204 4768 138256 4820
rect 164884 4768 164936 4820
rect 165712 4768 165764 4820
rect 527824 4768 527876 4820
rect 138940 4360 138992 4412
rect 143540 4360 143592 4412
rect 242900 4156 242952 4208
rect 244096 4156 244148 4208
rect 251180 4156 251232 4208
rect 252376 4156 252428 4208
rect 276020 4156 276072 4208
rect 276756 4156 276808 4208
rect 119896 4088 119948 4140
rect 124864 4088 124916 4140
rect 125876 4088 125928 4140
rect 134524 4088 134576 4140
rect 151544 4088 151596 4140
rect 325608 4088 325660 4140
rect 138664 4020 138716 4072
rect 145932 4020 145984 4072
rect 150532 4020 150584 4072
rect 328000 4020 328052 4072
rect 12348 3952 12400 4004
rect 126612 3952 126664 4004
rect 135812 3952 135864 4004
rect 141240 3952 141292 4004
rect 150900 3952 150952 4004
rect 331588 3952 331640 4004
rect 137744 3884 137796 3936
rect 144736 3884 144788 3936
rect 172152 3884 172204 3936
rect 356336 3884 356388 3936
rect 467104 3884 467156 3936
rect 534908 3884 534960 3936
rect 83280 3816 83332 3868
rect 131856 3816 131908 3868
rect 135536 3816 135588 3868
rect 138848 3816 138900 3868
rect 142988 3816 143040 3868
rect 151820 3816 151872 3868
rect 172060 3816 172112 3868
rect 303160 3816 303212 3868
rect 319444 3816 319496 3868
rect 583392 3816 583444 3868
rect 76196 3748 76248 3800
rect 129004 3748 129056 3800
rect 131764 3748 131816 3800
rect 135720 3748 135772 3800
rect 136824 3748 136876 3800
rect 69112 3680 69164 3732
rect 130660 3680 130712 3732
rect 135444 3680 135496 3732
rect 137652 3680 137704 3732
rect 140136 3748 140188 3800
rect 149520 3748 149572 3800
rect 152556 3748 152608 3800
rect 168380 3748 168432 3800
rect 178684 3748 178736 3800
rect 475752 3748 475804 3800
rect 154212 3680 154264 3732
rect 163964 3680 164016 3732
rect 491116 3680 491168 3732
rect 62028 3612 62080 3664
rect 122196 3612 122248 3664
rect 47860 3544 47912 3596
rect 127624 3612 127676 3664
rect 132960 3612 133012 3664
rect 135628 3612 135680 3664
rect 135904 3612 135956 3664
rect 140044 3612 140096 3664
rect 126980 3544 127032 3596
rect 130384 3544 130436 3596
rect 135352 3544 135404 3596
rect 136456 3544 136508 3596
rect 136732 3544 136784 3596
rect 155408 3612 155460 3664
rect 171876 3612 171928 3664
rect 501788 3612 501840 3664
rect 17040 3476 17092 3528
rect 126428 3476 126480 3528
rect 133788 3476 133840 3528
rect 147128 3544 147180 3596
rect 147220 3544 147272 3596
rect 167184 3544 167236 3596
rect 171784 3544 171836 3596
rect 515956 3544 516008 3596
rect 141516 3476 141568 3528
rect 166080 3476 166132 3528
rect 173164 3476 173216 3528
rect 93860 3408 93912 3460
rect 94780 3408 94832 3460
rect 142804 3408 142856 3460
rect 170772 3408 170824 3460
rect 173348 3408 173400 3460
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 150808 3340 150860 3392
rect 322112 3340 322164 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 506480 3340 506532 3392
rect 507308 3340 507360 3392
rect 533712 3408 533764 3460
rect 537208 3340 537260 3392
rect 144460 3272 144512 3324
rect 153016 3272 153068 3324
rect 173256 3272 173308 3324
rect 212172 3272 212224 3324
rect 211804 3204 211856 3256
rect 362316 3272 362368 3324
rect 307760 3204 307812 3256
rect 309048 3204 309100 3256
rect 316040 3204 316092 3256
rect 317328 3204 317380 3256
rect 390560 1232 390612 1284
rect 391848 1232 391900 1284
rect 30104 1096 30156 1148
rect 33232 1096 33284 1148
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3238 410544 3294 410553
rect 3238 410479 3240 410488
rect 3292 410479 3294 410488
rect 3240 410450 3292 410456
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3252 371278 3280 371311
rect 3240 371272 3292 371278
rect 3240 371214 3292 371220
rect 3238 358456 3294 358465
rect 3238 358391 3294 358400
rect 3252 357474 3280 358391
rect 3240 357468 3292 357474
rect 3240 357410 3292 357416
rect 3238 319288 3294 319297
rect 3238 319223 3294 319232
rect 3252 318850 3280 319223
rect 3240 318844 3292 318850
rect 3240 318786 3292 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292670 2820 293111
rect 2780 292664 2832 292670
rect 2780 292606 2832 292612
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 2870 228032 2926 228041
rect 2870 227967 2926 227976
rect 2884 227798 2912 227967
rect 2872 227792 2924 227798
rect 2872 227734 2924 227740
rect 3252 149734 3280 306167
rect 3344 231198 3372 423535
rect 3332 231192 3384 231198
rect 3332 231134 3384 231140
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 201920 3386 201929
rect 3330 201855 3332 201864
rect 3384 201855 3386 201864
rect 3332 201826 3384 201832
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 3240 149728 3292 149734
rect 3240 149670 3292 149676
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3332 135312 3384 135318
rect 3332 135254 3384 135260
rect 3240 133952 3292 133958
rect 3240 133894 3292 133900
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3252 97617 3280 133894
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3344 93854 3372 135254
rect 3160 93826 3372 93854
rect 3160 89714 3188 93826
rect 3068 89686 3188 89714
rect 3068 84862 3096 89686
rect 3148 85604 3200 85610
rect 3148 85546 3200 85552
rect 3056 84856 3108 84862
rect 3056 84798 3108 84804
rect 3160 80481 3188 85546
rect 3436 84946 3464 658135
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579698 3556 579935
rect 3516 579692 3568 579698
rect 3516 579634 3568 579640
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3528 85610 3556 553823
rect 3620 85610 3648 606047
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3516 85604 3568 85610
rect 3516 85546 3568 85552
rect 3608 85604 3660 85610
rect 3608 85546 3660 85552
rect 3712 85490 3740 449511
rect 3252 84918 3464 84946
rect 3528 85462 3740 85490
rect 3146 80472 3202 80481
rect 3146 80407 3202 80416
rect 3252 78985 3280 84918
rect 3332 84856 3384 84862
rect 3332 84798 3384 84804
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 1398 76528 1454 76537
rect 1398 76463 1454 76472
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 584 480 612 8910
rect 542 -960 654 480
rect 1412 354 1440 76463
rect 2778 75168 2834 75177
rect 2778 75103 2834 75112
rect 2792 16574 2820 75103
rect 3344 58585 3372 84798
rect 3528 81297 3556 85462
rect 3608 85400 3660 85406
rect 3608 85342 3660 85348
rect 3514 81288 3570 81297
rect 3514 81223 3570 81232
rect 3620 81138 3648 85342
rect 3804 85082 3832 501735
rect 4066 475688 4122 475697
rect 4066 475623 4122 475632
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 3882 345400 3938 345409
rect 3882 345335 3938 345344
rect 3436 81110 3648 81138
rect 3712 85054 3832 85082
rect 3436 79121 3464 81110
rect 3712 80054 3740 85054
rect 3896 84998 3924 345335
rect 3884 84992 3936 84998
rect 3884 84934 3936 84940
rect 3988 84810 4016 397423
rect 4080 231130 4108 475623
rect 4068 231124 4120 231130
rect 4068 231066 4120 231072
rect 4066 149832 4122 149841
rect 4066 149767 4122 149776
rect 4080 138718 4108 149767
rect 4816 140214 4844 683674
rect 4896 632120 4948 632126
rect 4896 632062 4948 632068
rect 4908 141642 4936 632062
rect 6184 527196 6236 527202
rect 6184 527138 6236 527144
rect 4988 462596 5040 462602
rect 4988 462538 5040 462544
rect 4896 141636 4948 141642
rect 4896 141578 4948 141584
rect 4804 140208 4856 140214
rect 4804 140150 4856 140156
rect 4068 138712 4120 138718
rect 4068 138654 4120 138660
rect 4068 136740 4120 136746
rect 4068 136682 4120 136688
rect 3620 80026 3740 80054
rect 3804 84782 4016 84810
rect 3620 79257 3648 80026
rect 3804 79393 3832 84782
rect 3884 84720 3936 84726
rect 3884 84662 3936 84668
rect 3974 84688 4030 84697
rect 3896 80617 3924 84662
rect 3974 84623 4030 84632
rect 3988 84250 4016 84623
rect 3976 84244 4028 84250
rect 3976 84186 4028 84192
rect 3882 80608 3938 80617
rect 3882 80543 3938 80552
rect 3790 79384 3846 79393
rect 3790 79319 3846 79328
rect 3606 79248 3662 79257
rect 3606 79183 3662 79192
rect 3422 79112 3478 79121
rect 3422 79047 3478 79056
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3436 32473 3464 32982
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 3436 6497 3464 23258
rect 4080 19417 4108 136682
rect 5000 124166 5028 462538
rect 5080 292664 5132 292670
rect 5080 292606 5132 292612
rect 4988 124160 5040 124166
rect 4988 124102 5040 124108
rect 5092 78878 5120 292606
rect 5172 240236 5224 240242
rect 5172 240178 5224 240184
rect 5184 79626 5212 240178
rect 6196 144362 6224 527138
rect 6184 144356 6236 144362
rect 6184 144298 6236 144304
rect 5172 79620 5224 79626
rect 5172 79562 5224 79568
rect 6932 79529 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 8944 410508 8996 410514
rect 8944 410450 8996 410456
rect 7564 201884 7616 201890
rect 7564 201826 7616 201832
rect 7576 131102 7604 201826
rect 7564 131096 7616 131102
rect 7564 131038 7616 131044
rect 8956 125594 8984 410450
rect 10336 140282 10364 579634
rect 10416 371272 10468 371278
rect 10416 371214 10468 371220
rect 10428 144430 10456 371214
rect 10416 144424 10468 144430
rect 10416 144366 10468 144372
rect 10324 140276 10376 140282
rect 10324 140218 10376 140224
rect 8944 125588 8996 125594
rect 8944 125530 8996 125536
rect 15856 118658 15884 670686
rect 19984 618316 20036 618322
rect 19984 618258 20036 618264
rect 19996 120086 20024 618258
rect 22744 357468 22796 357474
rect 22744 357410 22796 357416
rect 20076 266416 20128 266422
rect 20076 266358 20128 266364
rect 20088 162178 20116 266358
rect 20076 162172 20128 162178
rect 20076 162114 20128 162120
rect 22756 126954 22784 357410
rect 22836 253972 22888 253978
rect 22836 253914 22888 253920
rect 22848 129742 22876 253914
rect 22928 149728 22980 149734
rect 22928 149670 22980 149676
rect 22836 129736 22888 129742
rect 22836 129678 22888 129684
rect 22940 128314 22968 149670
rect 22928 128308 22980 128314
rect 22928 128250 22980 128256
rect 22744 126948 22796 126954
rect 22744 126890 22796 126896
rect 19984 120080 20036 120086
rect 19984 120022 20036 120028
rect 15844 118652 15896 118658
rect 15844 118594 15896 118600
rect 23492 117298 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 37924 565888 37976 565894
rect 37924 565830 37976 565836
rect 24124 514820 24176 514826
rect 24124 514762 24176 514768
rect 24136 122806 24164 514762
rect 33784 318844 33836 318850
rect 33784 318786 33836 318792
rect 33796 144498 33824 318786
rect 33784 144492 33836 144498
rect 33784 144434 33836 144440
rect 25504 138712 25556 138718
rect 25504 138654 25556 138660
rect 25516 132462 25544 138654
rect 25504 132456 25556 132462
rect 25504 132398 25556 132404
rect 24124 122800 24176 122806
rect 24124 122742 24176 122748
rect 37936 121446 37964 565830
rect 40052 141710 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 69664 396772 69716 396778
rect 69664 396714 69716 396720
rect 69676 385014 69704 396714
rect 68284 385008 68336 385014
rect 68284 384950 68336 384956
rect 69664 385008 69716 385014
rect 69664 384950 69716 384956
rect 59268 370524 59320 370530
rect 59268 370466 59320 370472
rect 59280 366382 59308 370466
rect 46940 366376 46992 366382
rect 46940 366318 46992 366324
rect 59268 366376 59320 366382
rect 59268 366318 59320 366324
rect 46952 361010 46980 366318
rect 45100 361004 45152 361010
rect 45100 360946 45152 360952
rect 46940 361004 46992 361010
rect 46940 360946 46992 360952
rect 44916 274712 44968 274718
rect 44916 274654 44968 274660
rect 44824 239828 44876 239834
rect 44824 239770 44876 239776
rect 44836 233034 44864 239770
rect 44824 233028 44876 233034
rect 44824 232970 44876 232976
rect 44928 220862 44956 274654
rect 45008 254312 45060 254318
rect 45008 254254 45060 254260
rect 44916 220856 44968 220862
rect 44916 220798 44968 220804
rect 45020 216646 45048 254254
rect 45112 217326 45140 360946
rect 68296 358834 68324 384950
rect 65432 358828 65484 358834
rect 65432 358770 65484 358776
rect 68284 358828 68336 358834
rect 68284 358770 68336 358776
rect 65444 358154 65472 358770
rect 64144 358148 64196 358154
rect 64144 358090 64196 358096
rect 65432 358148 65484 358154
rect 65432 358090 65484 358096
rect 63868 345704 63920 345710
rect 63868 345646 63920 345652
rect 63880 339250 63908 345646
rect 61384 339244 61436 339250
rect 61384 339186 61436 339192
rect 63868 339244 63920 339250
rect 63868 339186 63920 339192
rect 61396 314702 61424 339186
rect 62856 331900 62908 331906
rect 62856 331842 62908 331848
rect 62764 319456 62816 319462
rect 62764 319398 62816 319404
rect 61476 318436 61528 318442
rect 61476 318378 61528 318384
rect 58624 314696 58676 314702
rect 58624 314638 58676 314644
rect 61384 314696 61436 314702
rect 61384 314638 61436 314644
rect 53840 291848 53892 291854
rect 53840 291790 53892 291796
rect 53852 289882 53880 291790
rect 53840 289876 53892 289882
rect 53840 289818 53892 289824
rect 51816 289808 51868 289814
rect 51816 289750 51868 289756
rect 51828 280226 51856 289750
rect 57244 287700 57296 287706
rect 57244 287642 57296 287648
rect 55588 284300 55640 284306
rect 55588 284242 55640 284248
rect 55600 281178 55628 284242
rect 54208 281172 54260 281178
rect 54208 281114 54260 281120
rect 55588 281172 55640 281178
rect 55588 281114 55640 281120
rect 53288 280832 53340 280838
rect 53288 280774 53340 280780
rect 49700 280220 49752 280226
rect 49700 280162 49752 280168
rect 51816 280220 51868 280226
rect 51816 280162 51868 280168
rect 49712 278186 49740 280162
rect 53104 278860 53156 278866
rect 53104 278802 53156 278808
rect 48964 278180 49016 278186
rect 48964 278122 49016 278128
rect 49700 278180 49752 278186
rect 49700 278122 49752 278128
rect 46940 278044 46992 278050
rect 46940 277986 46992 277992
rect 46952 274718 46980 277986
rect 46940 274712 46992 274718
rect 46940 274654 46992 274660
rect 48320 266348 48372 266354
rect 48320 266290 48372 266296
rect 48332 262290 48360 266290
rect 48240 262262 48360 262290
rect 48240 259282 48268 262262
rect 45744 259276 45796 259282
rect 45744 259218 45796 259224
rect 48228 259276 48280 259282
rect 48228 259218 48280 259224
rect 45560 255332 45612 255338
rect 45560 255274 45612 255280
rect 45192 249824 45244 249830
rect 45192 249766 45244 249772
rect 45204 230518 45232 249766
rect 45284 239896 45336 239902
rect 45284 239838 45336 239844
rect 45296 231062 45324 239838
rect 45468 239760 45520 239766
rect 45468 239702 45520 239708
rect 45376 238808 45428 238814
rect 45376 238750 45428 238756
rect 45388 232354 45416 238750
rect 45480 232422 45508 239702
rect 45468 232416 45520 232422
rect 45468 232358 45520 232364
rect 45376 232348 45428 232354
rect 45376 232290 45428 232296
rect 45284 231056 45336 231062
rect 45284 230998 45336 231004
rect 45192 230512 45244 230518
rect 45192 230454 45244 230460
rect 45100 217320 45152 217326
rect 45100 217262 45152 217268
rect 45008 216640 45060 216646
rect 45008 216582 45060 216588
rect 45572 147014 45600 255274
rect 45652 240780 45704 240786
rect 45652 240722 45704 240728
rect 45664 238814 45692 240722
rect 45652 238808 45704 238814
rect 45652 238750 45704 238756
rect 45756 233170 45784 259218
rect 46940 258596 46992 258602
rect 46940 258538 46992 258544
rect 46952 255338 46980 258538
rect 48228 256828 48280 256834
rect 48228 256770 48280 256776
rect 46940 255332 46992 255338
rect 46940 255274 46992 255280
rect 48240 254318 48268 256770
rect 48228 254312 48280 254318
rect 48228 254254 48280 254260
rect 47584 254040 47636 254046
rect 47584 253982 47636 253988
rect 46940 253972 46992 253978
rect 46940 253914 46992 253920
rect 46952 249830 46980 253914
rect 46940 249824 46992 249830
rect 46940 249766 46992 249772
rect 47596 245682 47624 253982
rect 48976 253978 49004 278122
rect 53116 272066 53144 278802
rect 53196 274712 53248 274718
rect 53196 274654 53248 274660
rect 51724 272060 51776 272066
rect 51724 272002 51776 272008
rect 53104 272060 53156 272066
rect 53104 272002 53156 272008
rect 51080 270496 51132 270502
rect 51080 270438 51132 270444
rect 51092 266422 51120 270438
rect 51080 266416 51132 266422
rect 51080 266358 51132 266364
rect 51736 263634 51764 272002
rect 53208 267734 53236 274654
rect 53300 270502 53328 280774
rect 54220 278866 54248 281114
rect 54208 278860 54260 278866
rect 54208 278802 54260 278808
rect 54484 278792 54536 278798
rect 54484 278734 54536 278740
rect 53840 277364 53892 277370
rect 53840 277306 53892 277312
rect 53852 274718 53880 277306
rect 53840 274712 53892 274718
rect 53840 274654 53892 274660
rect 53288 270496 53340 270502
rect 53288 270438 53340 270444
rect 53116 267706 53236 267734
rect 49700 263628 49752 263634
rect 49700 263570 49752 263576
rect 51724 263628 51776 263634
rect 51724 263570 51776 263576
rect 49712 258602 49740 263570
rect 49700 258596 49752 258602
rect 49700 258538 49752 258544
rect 50436 256692 50488 256698
rect 50436 256634 50488 256640
rect 50448 254046 50476 256634
rect 50436 254040 50488 254046
rect 50436 253982 50488 253988
rect 48964 253972 49016 253978
rect 48964 253914 49016 253920
rect 49056 253972 49108 253978
rect 49056 253914 49108 253920
rect 46572 245676 46624 245682
rect 46572 245618 46624 245624
rect 47584 245676 47636 245682
rect 47584 245618 47636 245624
rect 45836 240576 45888 240582
rect 45836 240518 45888 240524
rect 45744 233164 45796 233170
rect 45744 233106 45796 233112
rect 45652 233028 45704 233034
rect 45652 232970 45704 232976
rect 45664 230382 45692 232970
rect 45848 232422 45876 240518
rect 46584 239902 46612 245618
rect 49068 244322 49096 253914
rect 53116 252618 53144 267706
rect 54496 266490 54524 278734
rect 57256 277438 57284 287642
rect 57980 282940 58032 282946
rect 57980 282882 58032 282888
rect 57992 280242 58020 282882
rect 57900 280214 58020 280242
rect 57900 278798 57928 280214
rect 57888 278792 57940 278798
rect 57888 278734 57940 278740
rect 58636 278050 58664 314638
rect 61488 311234 61516 318378
rect 60004 311228 60056 311234
rect 60004 311170 60056 311176
rect 61476 311228 61528 311234
rect 61476 311170 61528 311176
rect 60016 290426 60044 311170
rect 62776 299470 62804 319398
rect 62868 318442 62896 331842
rect 64156 319462 64184 358090
rect 64144 319456 64196 319462
rect 64144 319398 64196 319404
rect 62856 318436 62908 318442
rect 62856 318378 62908 318384
rect 71044 313336 71096 313342
rect 71044 313278 71096 313284
rect 71056 305046 71084 313278
rect 69664 305040 69716 305046
rect 69664 304982 69716 304988
rect 71044 305040 71096 305046
rect 71044 304982 71096 304988
rect 69676 302258 69704 304982
rect 68284 302252 68336 302258
rect 68284 302194 68336 302200
rect 69664 302252 69716 302258
rect 69664 302194 69716 302200
rect 60832 299464 60884 299470
rect 60832 299406 60884 299412
rect 62764 299464 62816 299470
rect 62764 299406 62816 299412
rect 60844 294030 60872 299406
rect 68296 294234 68324 302194
rect 66260 294228 66312 294234
rect 66260 294170 66312 294176
rect 68284 294228 68336 294234
rect 68284 294170 68336 294176
rect 60096 294024 60148 294030
rect 60096 293966 60148 293972
rect 60832 294024 60884 294030
rect 60832 293966 60884 293972
rect 58716 290420 58768 290426
rect 58716 290362 58768 290368
rect 60004 290420 60056 290426
rect 60004 290362 60056 290368
rect 58728 284374 58756 290362
rect 58716 284368 58768 284374
rect 58716 284310 58768 284316
rect 60108 282946 60136 293966
rect 66272 292670 66300 294170
rect 63500 292664 63552 292670
rect 63500 292606 63552 292612
rect 66260 292664 66312 292670
rect 66260 292606 66312 292612
rect 63512 291854 63540 292606
rect 63500 291848 63552 291854
rect 63500 291790 63552 291796
rect 71792 287706 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 84200 452124 84252 452130
rect 84200 452066 84252 452072
rect 84212 447846 84240 452066
rect 75184 447840 75236 447846
rect 75184 447782 75236 447788
rect 84200 447840 84252 447846
rect 84200 447782 84252 447788
rect 75196 392018 75224 447782
rect 75276 403640 75328 403646
rect 75276 403582 75328 403588
rect 72424 392012 72476 392018
rect 72424 391954 72476 391960
rect 75184 392012 75236 392018
rect 75184 391954 75236 391960
rect 72436 370530 72464 391954
rect 72424 370524 72476 370530
rect 72424 370466 72476 370472
rect 75288 353326 75316 403582
rect 86224 382288 86276 382294
rect 86224 382230 86276 382236
rect 86236 359038 86264 382230
rect 84844 359032 84896 359038
rect 84844 358974 84896 358980
rect 86224 359032 86276 359038
rect 86224 358974 86276 358980
rect 71872 353320 71924 353326
rect 71872 353262 71924 353268
rect 75276 353320 75328 353326
rect 75276 353262 75328 353268
rect 71884 345710 71912 353262
rect 84856 351966 84884 358974
rect 84844 351960 84896 351966
rect 84844 351902 84896 351908
rect 82360 351892 82412 351898
rect 82360 351834 82412 351840
rect 82372 349178 82400 351834
rect 80704 349172 80756 349178
rect 80704 349114 80756 349120
rect 82360 349172 82412 349178
rect 82360 349114 82412 349120
rect 71872 345704 71924 345710
rect 71872 345646 71924 345652
rect 80716 320210 80744 349114
rect 88352 331906 88380 702406
rect 93492 559564 93544 559570
rect 93492 559506 93544 559512
rect 93504 552566 93532 559506
rect 90364 552560 90416 552566
rect 90364 552502 90416 552508
rect 93492 552560 93544 552566
rect 93492 552502 93544 552508
rect 90376 452130 90404 552502
rect 90364 452124 90416 452130
rect 90364 452066 90416 452072
rect 103520 423292 103572 423298
rect 103520 423234 103572 423240
rect 103532 417722 103560 423234
rect 101404 417716 101456 417722
rect 101404 417658 101456 417664
rect 103520 417716 103572 417722
rect 103520 417658 103572 417664
rect 95332 407788 95384 407794
rect 95332 407730 95384 407736
rect 95344 403646 95372 407730
rect 101416 405754 101444 417658
rect 101404 405748 101456 405754
rect 101404 405690 101456 405696
rect 97448 405680 97500 405686
rect 97448 405622 97500 405628
rect 95332 403640 95384 403646
rect 95332 403582 95384 403588
rect 97460 401674 97488 405622
rect 96068 401668 96120 401674
rect 96068 401610 96120 401616
rect 97448 401668 97500 401674
rect 97448 401610 97500 401616
rect 96080 397866 96108 401610
rect 94504 397860 94556 397866
rect 94504 397802 94556 397808
rect 96068 397860 96120 397866
rect 96068 397802 96120 397808
rect 94516 390794 94544 397802
rect 92480 390788 92532 390794
rect 92480 390730 92532 390736
rect 94504 390788 94556 390794
rect 94504 390730 94556 390736
rect 92492 385762 92520 390730
rect 90088 385756 90140 385762
rect 90088 385698 90140 385704
rect 92480 385756 92532 385762
rect 92480 385698 92532 385704
rect 90100 382294 90128 385698
rect 90088 382288 90140 382294
rect 90088 382230 90140 382236
rect 88340 331900 88392 331906
rect 88340 331842 88392 331848
rect 79508 320204 79560 320210
rect 79508 320146 79560 320152
rect 80704 320204 80756 320210
rect 80704 320146 80756 320152
rect 79520 318374 79548 320146
rect 78128 318368 78180 318374
rect 78128 318310 78180 318316
rect 79508 318368 79560 318374
rect 79508 318310 79560 318316
rect 78140 315314 78168 318310
rect 104912 315314 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136364 627904 136416 627910
rect 136364 627846 136416 627852
rect 136376 620362 136404 627846
rect 134524 620356 134576 620362
rect 134524 620298 134576 620304
rect 136364 620356 136416 620362
rect 136364 620298 136416 620304
rect 134536 608802 134564 620298
rect 126244 608796 126296 608802
rect 126244 608738 126296 608744
rect 134524 608796 134576 608802
rect 134524 608738 134576 608744
rect 126256 591326 126284 608738
rect 133144 592068 133196 592074
rect 133144 592010 133196 592016
rect 120724 591320 120776 591326
rect 120724 591262 120776 591268
rect 126244 591320 126296 591326
rect 126244 591262 126296 591268
rect 120736 585206 120764 591262
rect 119344 585200 119396 585206
rect 119344 585142 119396 585148
rect 120724 585200 120776 585206
rect 120724 585142 120776 585148
rect 119356 553450 119384 585142
rect 133156 578270 133184 592010
rect 129740 578264 129792 578270
rect 129740 578206 129792 578212
rect 133144 578264 133196 578270
rect 133144 578206 133196 578212
rect 129752 570654 129780 578206
rect 120724 570648 120776 570654
rect 120724 570590 120776 570596
rect 129740 570648 129792 570654
rect 129740 570590 129792 570596
rect 120736 559570 120764 570590
rect 120724 559564 120776 559570
rect 120724 559506 120776 559512
rect 117964 553444 118016 553450
rect 117964 553386 118016 553392
rect 119344 553444 119396 553450
rect 119344 553386 119396 553392
rect 117976 536858 118004 553386
rect 116584 536852 116636 536858
rect 116584 536794 116636 536800
rect 117964 536852 118016 536858
rect 117964 536794 118016 536800
rect 116596 534138 116624 536794
rect 115204 534132 115256 534138
rect 115204 534074 115256 534080
rect 116584 534132 116636 534138
rect 116584 534074 116636 534080
rect 115216 525842 115244 534074
rect 113824 525836 113876 525842
rect 113824 525778 113876 525784
rect 115204 525836 115256 525842
rect 115204 525778 115256 525784
rect 113836 481710 113864 525778
rect 112536 481704 112588 481710
rect 112536 481646 112588 481652
rect 113824 481704 113876 481710
rect 113824 481646 113876 481652
rect 112548 476134 112576 481646
rect 111064 476128 111116 476134
rect 111064 476070 111116 476076
rect 112536 476128 112588 476134
rect 112536 476070 112588 476076
rect 111076 459610 111104 476070
rect 109684 459604 109736 459610
rect 109684 459546 109736 459552
rect 111064 459604 111116 459610
rect 111064 459546 111116 459552
rect 109696 430642 109724 459546
rect 134708 431248 134760 431254
rect 134708 431190 134760 431196
rect 107660 430636 107712 430642
rect 107660 430578 107712 430584
rect 109684 430636 109736 430642
rect 109684 430578 109736 430584
rect 107672 427174 107700 430578
rect 106188 427168 106240 427174
rect 106188 427110 106240 427116
rect 107660 427168 107712 427174
rect 107660 427110 107712 427116
rect 106200 423298 106228 427110
rect 106188 423292 106240 423298
rect 106188 423234 106240 423240
rect 134720 422346 134748 431190
rect 131764 422340 131816 422346
rect 131764 422282 131816 422288
rect 134708 422340 134760 422346
rect 134708 422282 134760 422288
rect 131776 413302 131804 422282
rect 113180 413296 113232 413302
rect 113180 413238 113232 413244
rect 131764 413296 131816 413302
rect 131764 413238 131816 413244
rect 113192 407794 113220 413238
rect 113180 407788 113232 407794
rect 113180 407730 113232 407736
rect 136652 396778 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 699718 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 150440 699712 150492 699718
rect 150440 699654 150492 699660
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 150452 693530 150480 699654
rect 149796 693524 149848 693530
rect 149796 693466 149848 693472
rect 150440 693524 150492 693530
rect 150440 693466 150492 693472
rect 149808 687546 149836 693466
rect 148324 687540 148376 687546
rect 148324 687482 148376 687488
rect 149796 687540 149848 687546
rect 149796 687482 149848 687488
rect 148336 679046 148364 687482
rect 148324 679040 148376 679046
rect 148324 678982 148376 678988
rect 144184 678972 144236 678978
rect 144184 678914 144236 678920
rect 144196 662454 144224 678914
rect 167000 671356 167052 671362
rect 167000 671298 167052 671304
rect 167012 667214 167040 671298
rect 160744 667208 160796 667214
rect 160744 667150 160796 667156
rect 167000 667208 167052 667214
rect 167000 667150 167052 667156
rect 141424 662448 141476 662454
rect 141424 662390 141476 662396
rect 144184 662448 144236 662454
rect 144184 662390 144236 662396
rect 141436 638246 141464 662390
rect 160756 661094 160784 667150
rect 153844 661088 153896 661094
rect 153844 661030 153896 661036
rect 160744 661088 160796 661094
rect 160744 661030 160796 661036
rect 153856 652050 153884 661030
rect 146944 652044 146996 652050
rect 146944 651986 146996 651992
rect 153844 652044 153896 652050
rect 153844 651986 153896 651992
rect 146956 641782 146984 651986
rect 144184 641776 144236 641782
rect 144184 641718 144236 641724
rect 146944 641776 146996 641782
rect 146944 641718 146996 641724
rect 140044 638240 140096 638246
rect 140044 638182 140096 638188
rect 141424 638240 141476 638246
rect 141424 638182 141476 638188
rect 140056 627978 140084 638182
rect 140044 627972 140096 627978
rect 140044 627914 140096 627920
rect 144196 597582 144224 641718
rect 137744 597576 137796 597582
rect 137744 597518 137796 597524
rect 144184 597576 144236 597582
rect 144184 597518 144236 597524
rect 137756 592074 137784 597518
rect 137744 592068 137796 592074
rect 137744 592010 137796 592016
rect 167000 437436 167052 437442
rect 167000 437378 167052 437384
rect 151084 436756 151136 436762
rect 151084 436698 151136 436704
rect 151096 431254 151124 436698
rect 167012 434738 167040 437378
rect 166920 434710 167040 434738
rect 166920 433362 166948 434710
rect 166908 433356 166960 433362
rect 166908 433298 166960 433304
rect 163596 433288 163648 433294
rect 163596 433230 163648 433236
rect 151084 431248 151136 431254
rect 151084 431190 151136 431196
rect 163504 425740 163556 425746
rect 163504 425682 163556 425688
rect 160744 414044 160796 414050
rect 160744 413986 160796 413992
rect 148324 402280 148376 402286
rect 148324 402222 148376 402228
rect 136640 396772 136692 396778
rect 136640 396714 136692 396720
rect 148336 353326 148364 402222
rect 160756 366790 160784 413986
rect 163516 407114 163544 425682
rect 163608 414050 163636 433230
rect 163596 414044 163648 414050
rect 163596 413986 163648 413992
rect 160836 407108 160888 407114
rect 160836 407050 160888 407056
rect 163504 407108 163556 407114
rect 163504 407050 163556 407056
rect 160848 402286 160876 407050
rect 160836 402280 160888 402286
rect 160836 402222 160888 402228
rect 159364 366784 159416 366790
rect 159364 366726 159416 366732
rect 160744 366784 160796 366790
rect 160744 366726 160796 366732
rect 159376 356046 159404 366726
rect 157984 356040 158036 356046
rect 157984 355982 158036 355988
rect 159364 356040 159416 356046
rect 159364 355982 159416 355988
rect 145564 353320 145616 353326
rect 145564 353262 145616 353268
rect 148324 353320 148376 353326
rect 148324 353262 148376 353268
rect 145576 337414 145604 353262
rect 140412 337408 140464 337414
rect 140412 337350 140464 337356
rect 145564 337408 145616 337414
rect 145564 337350 145616 337356
rect 140424 328914 140452 337350
rect 157996 332654 158024 355982
rect 156696 332648 156748 332654
rect 156696 332590 156748 332596
rect 157984 332648 158036 332654
rect 157984 332590 158036 332596
rect 135904 328908 135956 328914
rect 135904 328850 135956 328856
rect 140412 328908 140464 328914
rect 140412 328850 140464 328856
rect 73160 315308 73212 315314
rect 73160 315250 73212 315256
rect 78128 315308 78180 315314
rect 78128 315250 78180 315256
rect 84844 315308 84896 315314
rect 84844 315250 84896 315256
rect 104900 315308 104952 315314
rect 104900 315250 104952 315256
rect 73172 313342 73200 315250
rect 73160 313336 73212 313342
rect 73160 313278 73212 313284
rect 71780 287700 71832 287706
rect 71780 287642 71832 287648
rect 82820 284980 82872 284986
rect 82820 284922 82872 284928
rect 82084 284300 82136 284306
rect 82084 284242 82136 284248
rect 60096 282940 60148 282946
rect 60096 282882 60148 282888
rect 66904 282192 66956 282198
rect 66904 282134 66956 282140
rect 58624 278044 58676 278050
rect 58624 277986 58676 277992
rect 57244 277432 57296 277438
rect 57244 277374 57296 277380
rect 55864 276684 55916 276690
rect 55864 276626 55916 276632
rect 53196 266484 53248 266490
rect 53196 266426 53248 266432
rect 54484 266484 54536 266490
rect 54484 266426 54536 266432
rect 53208 253978 53236 266426
rect 55876 266422 55904 276626
rect 66916 275126 66944 282134
rect 82096 276690 82124 284242
rect 82832 282198 82860 284922
rect 84856 284374 84884 315250
rect 135916 308446 135944 328850
rect 156708 328098 156736 332590
rect 155224 328092 155276 328098
rect 155224 328034 155276 328040
rect 156696 328092 156748 328098
rect 156696 328034 156748 328040
rect 155236 318782 155264 328034
rect 153844 318776 153896 318782
rect 153844 318718 153896 318724
rect 155224 318776 155276 318782
rect 155224 318718 155276 318724
rect 102784 308440 102836 308446
rect 102784 308382 102836 308388
rect 135904 308440 135956 308446
rect 135904 308382 135956 308388
rect 102796 297430 102824 308382
rect 153856 307834 153884 318718
rect 153844 307828 153896 307834
rect 153844 307770 153896 307776
rect 151084 307760 151136 307766
rect 151084 307702 151136 307708
rect 97724 297424 97776 297430
rect 97724 297366 97776 297372
rect 102784 297424 102836 297430
rect 102784 297366 102836 297372
rect 97736 294642 97764 297366
rect 87604 294636 87656 294642
rect 87604 294578 87656 294584
rect 97724 294636 97776 294642
rect 97724 294578 97776 294584
rect 87616 284986 87644 294578
rect 87604 284980 87656 284986
rect 87604 284922 87656 284928
rect 84844 284368 84896 284374
rect 84844 284310 84896 284316
rect 82820 282192 82872 282198
rect 82820 282134 82872 282140
rect 151096 281314 151124 307702
rect 148324 281308 148376 281314
rect 148324 281250 148376 281256
rect 151084 281308 151136 281314
rect 151084 281250 151136 281256
rect 82084 276684 82136 276690
rect 82084 276626 82136 276632
rect 63500 275120 63552 275126
rect 63500 275062 63552 275068
rect 66904 275120 66956 275126
rect 66904 275062 66956 275068
rect 63512 268666 63540 275062
rect 60556 268660 60608 268666
rect 60556 268602 60608 268608
rect 63500 268660 63552 268666
rect 63500 268602 63552 268608
rect 54208 266416 54260 266422
rect 54208 266358 54260 266364
rect 55864 266416 55916 266422
rect 55864 266358 55916 266364
rect 54220 263634 54248 266358
rect 53288 263628 53340 263634
rect 53288 263570 53340 263576
rect 54208 263628 54260 263634
rect 54208 263570 54260 263576
rect 53300 256766 53328 263570
rect 60568 262886 60596 268602
rect 148336 262954 148364 281250
rect 169772 280838 169800 702406
rect 202800 699718 202828 703520
rect 195980 699712 196032 699718
rect 195980 699654 196032 699660
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 195992 694822 196020 699654
rect 189080 694816 189132 694822
rect 189080 694758 189132 694764
rect 195980 694816 196032 694822
rect 195980 694758 196032 694764
rect 189092 688702 189120 694758
rect 181444 688696 181496 688702
rect 181444 688638 181496 688644
rect 189080 688696 189132 688702
rect 189080 688638 189132 688644
rect 181456 671362 181484 688638
rect 218072 687954 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 699718 235212 703520
rect 231860 699712 231912 699718
rect 231860 699654 231912 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 231872 695298 231900 699654
rect 229744 695292 229796 695298
rect 229744 695234 229796 695240
rect 231860 695292 231912 695298
rect 231860 695234 231912 695240
rect 206284 687948 206336 687954
rect 206284 687890 206336 687896
rect 218060 687948 218112 687954
rect 218060 687890 218112 687896
rect 206296 681766 206324 687890
rect 229756 685166 229784 695234
rect 267660 694278 267688 703520
rect 283852 698358 283880 703520
rect 281540 698352 281592 698358
rect 281540 698294 281592 698300
rect 283840 698352 283892 698358
rect 283840 698294 283892 698300
rect 281552 695026 281580 698294
rect 300136 698154 300164 703520
rect 332520 699854 332548 703520
rect 332508 699848 332560 699854
rect 332508 699790 332560 699796
rect 334624 699848 334676 699854
rect 334624 699790 334676 699796
rect 300124 698148 300176 698154
rect 300124 698090 300176 698096
rect 302884 698148 302936 698154
rect 302884 698090 302936 698096
rect 280804 695020 280856 695026
rect 280804 694962 280856 694968
rect 281540 695020 281592 695026
rect 281540 694962 281592 694968
rect 258080 694272 258132 694278
rect 258080 694214 258132 694220
rect 267648 694272 267700 694278
rect 267648 694214 267700 694220
rect 258092 689314 258120 694214
rect 247684 689308 247736 689314
rect 247684 689250 247736 689256
rect 258080 689308 258132 689314
rect 258080 689250 258132 689256
rect 221464 685160 221516 685166
rect 221464 685102 221516 685108
rect 229744 685160 229796 685166
rect 229744 685102 229796 685108
rect 204260 681760 204312 681766
rect 204260 681702 204312 681708
rect 206284 681760 206336 681766
rect 206284 681702 206336 681708
rect 204272 677074 204300 681702
rect 202144 677068 202196 677074
rect 202144 677010 202196 677016
rect 204260 677068 204312 677074
rect 204260 677010 204312 677016
rect 181444 671356 181496 671362
rect 181444 671298 181496 671304
rect 202156 666398 202184 677010
rect 221476 668642 221504 685102
rect 215944 668636 215996 668642
rect 215944 668578 215996 668584
rect 221464 668636 221516 668642
rect 221464 668578 221516 668584
rect 200120 666392 200172 666398
rect 200120 666334 200172 666340
rect 202144 666392 202196 666398
rect 202144 666334 202196 666340
rect 200132 659258 200160 666334
rect 195152 659252 195204 659258
rect 195152 659194 195204 659200
rect 200120 659252 200172 659258
rect 200120 659194 200172 659200
rect 195164 654838 195192 659194
rect 185584 654832 185636 654838
rect 185584 654774 185636 654780
rect 195152 654832 195204 654838
rect 195152 654774 195204 654780
rect 185596 632126 185624 654774
rect 215956 647902 215984 668578
rect 247696 658986 247724 689250
rect 280816 665174 280844 694962
rect 302896 692102 302924 698090
rect 302884 692096 302936 692102
rect 302884 692038 302936 692044
rect 313924 692096 313976 692102
rect 313924 692038 313976 692044
rect 313936 682446 313964 692038
rect 334636 686526 334664 699790
rect 348804 699718 348832 703520
rect 364996 700330 365024 703520
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 374644 700324 374696 700330
rect 374644 700266 374696 700272
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 350540 699712 350592 699718
rect 350540 699654 350592 699660
rect 350552 698086 350580 699654
rect 350540 698080 350592 698086
rect 350540 698022 350592 698028
rect 353944 698080 353996 698086
rect 353944 698022 353996 698028
rect 334624 686520 334676 686526
rect 334624 686462 334676 686468
rect 349804 686520 349856 686526
rect 349804 686462 349856 686468
rect 313924 682440 313976 682446
rect 313924 682382 313976 682388
rect 333244 682440 333296 682446
rect 333244 682382 333296 682388
rect 279424 665168 279476 665174
rect 279424 665110 279476 665116
rect 280804 665168 280856 665174
rect 280804 665110 280856 665116
rect 241980 658980 242032 658986
rect 241980 658922 242032 658928
rect 247684 658980 247736 658986
rect 247684 658922 247736 658928
rect 241992 656198 242020 658922
rect 235264 656192 235316 656198
rect 235264 656134 235316 656140
rect 241980 656192 242032 656198
rect 241980 656134 242032 656140
rect 203524 647896 203576 647902
rect 203524 647838 203576 647844
rect 215944 647896 215996 647902
rect 215944 647838 215996 647844
rect 203536 635526 203564 647838
rect 235276 639470 235304 656134
rect 279436 655586 279464 665110
rect 274640 655580 274692 655586
rect 274640 655522 274692 655528
rect 279424 655580 279476 655586
rect 279424 655522 279476 655528
rect 274652 652798 274680 655522
rect 273904 652792 273956 652798
rect 273904 652734 273956 652740
rect 274640 652792 274692 652798
rect 274640 652734 274692 652740
rect 232504 639464 232556 639470
rect 232504 639406 232556 639412
rect 235264 639464 235316 639470
rect 235264 639406 235316 639412
rect 196624 635520 196676 635526
rect 196624 635462 196676 635468
rect 203524 635520 203576 635526
rect 203524 635462 203576 635468
rect 184204 632120 184256 632126
rect 184204 632062 184256 632068
rect 185584 632120 185636 632126
rect 185584 632062 185636 632068
rect 184216 603158 184244 632062
rect 182824 603152 182876 603158
rect 182824 603094 182876 603100
rect 184204 603152 184256 603158
rect 184204 603094 184256 603100
rect 182836 578202 182864 603094
rect 181444 578196 181496 578202
rect 181444 578138 181496 578144
rect 182824 578196 182876 578202
rect 182824 578138 182876 578144
rect 181456 524482 181484 578138
rect 196636 554810 196664 635462
rect 232516 590374 232544 639406
rect 273916 632126 273944 652734
rect 333256 643754 333284 682382
rect 349816 658238 349844 686462
rect 353956 683806 353984 698022
rect 374656 691150 374684 700266
rect 374644 691144 374696 691150
rect 374644 691086 374696 691092
rect 377404 691144 377456 691150
rect 377404 691086 377456 691092
rect 353944 683800 353996 683806
rect 353944 683742 353996 683748
rect 358360 683800 358412 683806
rect 358360 683742 358412 683748
rect 358372 678502 358400 683742
rect 358360 678496 358412 678502
rect 358360 678438 358412 678444
rect 360844 678496 360896 678502
rect 360844 678438 360896 678444
rect 360856 668642 360884 678438
rect 377416 678298 377444 691086
rect 377404 678292 377456 678298
rect 377404 678234 377456 678240
rect 396448 678292 396500 678298
rect 396448 678234 396500 678240
rect 360844 668636 360896 668642
rect 360844 668578 360896 668584
rect 363604 668636 363656 668642
rect 363604 668578 363656 668584
rect 363616 663066 363644 668578
rect 363604 663060 363656 663066
rect 363604 663002 363656 663008
rect 369124 663060 369176 663066
rect 369124 663002 369176 663008
rect 369136 660346 369164 663002
rect 369124 660340 369176 660346
rect 369124 660282 369176 660288
rect 387340 660340 387392 660346
rect 387340 660282 387392 660288
rect 387352 658238 387380 660282
rect 349804 658232 349856 658238
rect 349804 658174 349856 658180
rect 355784 658232 355836 658238
rect 355784 658174 355836 658180
rect 387340 658232 387392 658238
rect 387340 658174 387392 658180
rect 393964 658232 394016 658238
rect 393964 658174 394016 658180
rect 355796 655518 355824 658174
rect 355784 655512 355836 655518
rect 355784 655454 355836 655460
rect 358728 655512 358780 655518
rect 358728 655454 358780 655460
rect 358740 650690 358768 655454
rect 358728 650684 358780 650690
rect 358728 650626 358780 650632
rect 369124 650684 369176 650690
rect 369124 650626 369176 650632
rect 333244 643748 333296 643754
rect 333244 643690 333296 643696
rect 353944 643748 353996 643754
rect 353944 643690 353996 643696
rect 272616 632120 272668 632126
rect 272616 632062 272668 632068
rect 273904 632120 273956 632126
rect 273904 632062 273956 632068
rect 272628 629746 272656 632062
rect 271144 629740 271196 629746
rect 271144 629682 271196 629688
rect 272616 629740 272668 629746
rect 272616 629682 272668 629688
rect 271156 616826 271184 629682
rect 353956 625870 353984 643690
rect 369136 640558 369164 650626
rect 393976 649942 394004 658174
rect 393964 649936 394016 649942
rect 393964 649878 394016 649884
rect 395344 649936 395396 649942
rect 395344 649878 395396 649884
rect 395356 647222 395384 649878
rect 395344 647216 395396 647222
rect 395344 647158 395396 647164
rect 369124 640552 369176 640558
rect 369124 640494 369176 640500
rect 371884 640552 371936 640558
rect 371884 640494 371936 640500
rect 353944 625864 353996 625870
rect 353944 625806 353996 625812
rect 269396 616820 269448 616826
rect 269396 616762 269448 616768
rect 271144 616820 271196 616826
rect 271144 616762 271196 616768
rect 269408 608802 269436 616762
rect 268384 608796 268436 608802
rect 268384 608738 268436 608744
rect 269396 608796 269448 608802
rect 269396 608738 269448 608744
rect 268396 593570 268424 608738
rect 264244 593564 264296 593570
rect 264244 593506 264296 593512
rect 268384 593564 268436 593570
rect 268384 593506 268436 593512
rect 229744 590368 229796 590374
rect 229744 590310 229796 590316
rect 232504 590368 232556 590374
rect 232504 590310 232556 590316
rect 229756 581670 229784 590310
rect 264256 585206 264284 593506
rect 371896 591326 371924 640494
rect 395344 625864 395396 625870
rect 395344 625806 395396 625812
rect 371884 591320 371936 591326
rect 371884 591262 371936 591268
rect 384304 591320 384356 591326
rect 384304 591262 384356 591268
rect 262864 585200 262916 585206
rect 262864 585142 262916 585148
rect 264244 585200 264296 585206
rect 264244 585142 264296 585148
rect 207664 581664 207716 581670
rect 207664 581606 207716 581612
rect 229744 581664 229796 581670
rect 229744 581606 229796 581612
rect 193864 554804 193916 554810
rect 193864 554746 193916 554752
rect 196624 554804 196676 554810
rect 196624 554746 196676 554752
rect 181444 524476 181496 524482
rect 181444 524418 181496 524424
rect 177304 524408 177356 524414
rect 177304 524350 177356 524356
rect 177316 505170 177344 524350
rect 193876 520266 193904 554746
rect 207676 545766 207704 581606
rect 262876 570654 262904 585142
rect 384316 583574 384344 591262
rect 384304 583568 384356 583574
rect 384304 583510 384356 583516
rect 390560 583568 390612 583574
rect 390560 583510 390612 583516
rect 390572 576910 390600 583510
rect 390560 576904 390612 576910
rect 390560 576846 390612 576852
rect 393964 576904 394016 576910
rect 393964 576846 394016 576852
rect 261484 570648 261536 570654
rect 261484 570590 261536 570596
rect 262864 570648 262916 570654
rect 262864 570590 262916 570596
rect 261496 552158 261524 570590
rect 260196 552152 260248 552158
rect 260196 552094 260248 552100
rect 261484 552152 261536 552158
rect 261484 552094 261536 552100
rect 260208 550050 260236 552094
rect 258816 550044 258868 550050
rect 258816 549986 258868 549992
rect 260196 550044 260248 550050
rect 260196 549986 260248 549992
rect 198004 545760 198056 545766
rect 198004 545702 198056 545708
rect 207664 545760 207716 545766
rect 207664 545702 207716 545708
rect 191104 520260 191156 520266
rect 191104 520202 191156 520208
rect 193864 520260 193916 520266
rect 193864 520202 193916 520208
rect 173164 505164 173216 505170
rect 173164 505106 173216 505112
rect 177304 505164 177356 505170
rect 177304 505106 177356 505112
rect 173176 473074 173204 505106
rect 171784 473068 171836 473074
rect 171784 473010 171836 473016
rect 173164 473068 173216 473074
rect 173164 473010 173216 473016
rect 171796 447098 171824 473010
rect 189080 470620 189132 470626
rect 189080 470562 189132 470568
rect 189092 466478 189120 470562
rect 182824 466472 182876 466478
rect 182824 466414 182876 466420
rect 189080 466472 189132 466478
rect 189080 466414 189132 466420
rect 182836 459610 182864 466414
rect 179420 459604 179472 459610
rect 179420 459546 179472 459552
rect 182824 459604 182876 459610
rect 182824 459546 182876 459552
rect 179432 452606 179460 459546
rect 177304 452600 177356 452606
rect 177304 452542 177356 452548
rect 179420 452600 179472 452606
rect 179420 452542 179472 452548
rect 170404 447092 170456 447098
rect 170404 447034 170456 447040
rect 171784 447092 171836 447098
rect 171784 447034 171836 447040
rect 170416 437510 170444 447034
rect 170404 437504 170456 437510
rect 170404 437446 170456 437452
rect 177316 436762 177344 452542
rect 177304 436756 177356 436762
rect 177304 436698 177356 436704
rect 191116 429894 191144 520202
rect 198016 504422 198044 545702
rect 258828 542026 258856 549986
rect 256700 542020 256752 542026
rect 256700 541962 256752 541968
rect 258816 542020 258868 542026
rect 258816 541962 258868 541968
rect 256712 538898 256740 541962
rect 255964 538892 256016 538898
rect 255964 538834 256016 538840
rect 256700 538892 256752 538898
rect 256700 538834 256752 538840
rect 255976 511834 256004 538834
rect 393976 536450 394004 576846
rect 393964 536444 394016 536450
rect 393964 536386 394016 536392
rect 253940 511828 253992 511834
rect 253940 511770 253992 511776
rect 255964 511828 256016 511834
rect 255964 511770 256016 511776
rect 253952 506530 253980 511770
rect 251824 506524 251876 506530
rect 251824 506466 251876 506472
rect 253940 506524 253992 506530
rect 253940 506466 253992 506472
rect 195244 504416 195296 504422
rect 195244 504358 195296 504364
rect 198004 504416 198056 504422
rect 198004 504358 198056 504364
rect 195256 490074 195284 504358
rect 192484 490068 192536 490074
rect 192484 490010 192536 490016
rect 195244 490068 195296 490074
rect 195244 490010 195296 490016
rect 192496 470626 192524 490010
rect 192484 470620 192536 470626
rect 192484 470562 192536 470568
rect 251836 466478 251864 506466
rect 250168 466472 250220 466478
rect 250168 466414 250220 466420
rect 251824 466472 251876 466478
rect 251824 466414 251876 466420
rect 250180 463010 250208 466414
rect 248420 463004 248472 463010
rect 248420 462946 248472 462952
rect 250168 463004 250220 463010
rect 250168 462946 250220 462952
rect 248432 459610 248460 462946
rect 245752 459604 245804 459610
rect 245752 459546 245804 459552
rect 248420 459604 248472 459610
rect 248420 459546 248472 459552
rect 245764 455462 245792 459546
rect 244924 455456 244976 455462
rect 244924 455398 244976 455404
rect 245752 455456 245804 455462
rect 245752 455398 245804 455404
rect 171508 429888 171560 429894
rect 171508 429830 171560 429836
rect 191104 429888 191156 429894
rect 191104 429830 191156 429836
rect 171520 425746 171548 429830
rect 171508 425740 171560 425746
rect 171508 425682 171560 425688
rect 244936 416770 244964 455398
rect 243544 416764 243596 416770
rect 243544 416706 243596 416712
rect 244924 416764 244976 416770
rect 244924 416706 244976 416712
rect 243556 403646 243584 416706
rect 236644 403640 236696 403646
rect 236644 403582 236696 403588
rect 243544 403640 243596 403646
rect 243544 403582 243596 403588
rect 236656 396030 236684 403582
rect 233884 396024 233936 396030
rect 233884 395966 233936 395972
rect 236644 396024 236696 396030
rect 236644 395966 236696 395972
rect 233896 349858 233924 395966
rect 228364 349852 228416 349858
rect 228364 349794 228416 349800
rect 233884 349852 233936 349858
rect 233884 349794 233936 349800
rect 228376 338094 228404 349794
rect 225604 338088 225656 338094
rect 225604 338030 225656 338036
rect 228364 338088 228416 338094
rect 228364 338030 228416 338036
rect 225616 317422 225644 338030
rect 224224 317416 224276 317422
rect 224224 317358 224276 317364
rect 225604 317416 225656 317422
rect 225604 317358 225656 317364
rect 224236 303686 224264 317358
rect 224224 303680 224276 303686
rect 224224 303622 224276 303628
rect 220820 303612 220872 303618
rect 220820 303554 220872 303560
rect 220832 301170 220860 303554
rect 220084 301164 220136 301170
rect 220084 301106 220136 301112
rect 220820 301164 220872 301170
rect 220820 301106 220872 301112
rect 220096 291242 220124 301106
rect 220084 291236 220136 291242
rect 220084 291178 220136 291184
rect 213828 291168 213880 291174
rect 213828 291110 213880 291116
rect 213840 288930 213868 291110
rect 211160 288924 211212 288930
rect 211160 288866 211212 288872
rect 213828 288924 213880 288930
rect 213828 288866 213880 288872
rect 211172 284034 211200 288866
rect 207020 284028 207072 284034
rect 207020 283970 207072 283976
rect 211160 284028 211212 284034
rect 211160 283970 211212 283976
rect 169760 280832 169812 280838
rect 169760 280774 169812 280780
rect 207032 278322 207060 283970
rect 204168 278316 204220 278322
rect 204168 278258 204220 278264
rect 207020 278316 207072 278322
rect 207020 278258 207072 278264
rect 204180 274718 204208 278258
rect 201500 274712 201552 274718
rect 201500 274654 201552 274660
rect 204168 274712 204220 274718
rect 204168 274654 204220 274660
rect 201512 270978 201540 274654
rect 200764 270972 200816 270978
rect 200764 270914 200816 270920
rect 201500 270972 201552 270978
rect 201500 270914 201552 270920
rect 200776 266422 200804 270914
rect 198004 266416 198056 266422
rect 198004 266358 198056 266364
rect 200764 266416 200816 266422
rect 200764 266358 200816 266364
rect 146944 262948 146996 262954
rect 146944 262890 146996 262896
rect 148324 262948 148376 262954
rect 148324 262890 148376 262896
rect 53380 262880 53432 262886
rect 53380 262822 53432 262828
rect 60556 262880 60608 262886
rect 60556 262822 60608 262828
rect 53392 256834 53420 262822
rect 53380 256828 53432 256834
rect 53380 256770 53432 256776
rect 53288 256760 53340 256766
rect 53288 256702 53340 256708
rect 146956 253978 146984 262890
rect 53196 253972 53248 253978
rect 53196 253914 53248 253920
rect 144276 253972 144328 253978
rect 144276 253914 144328 253920
rect 146944 253972 146996 253978
rect 146944 253914 146996 253920
rect 144288 252890 144316 253914
rect 135904 252884 135956 252890
rect 135904 252826 135956 252832
rect 144276 252884 144328 252890
rect 144276 252826 144328 252832
rect 51816 252612 51868 252618
rect 51816 252554 51868 252560
rect 53104 252612 53156 252618
rect 53104 252554 53156 252560
rect 51828 250714 51856 252554
rect 50344 250708 50396 250714
rect 50344 250650 50396 250656
rect 51816 250708 51868 250714
rect 51816 250650 51868 250656
rect 46940 244316 46992 244322
rect 46940 244258 46992 244264
rect 49056 244316 49108 244322
rect 49056 244258 49108 244264
rect 46952 241618 46980 244258
rect 46768 241590 46980 241618
rect 46572 239896 46624 239902
rect 46572 239838 46624 239844
rect 46768 239766 46796 241590
rect 46848 240848 46900 240854
rect 46848 240790 46900 240796
rect 46860 239834 46888 240790
rect 50356 240582 50384 250650
rect 135916 243098 135944 252826
rect 198016 245682 198044 266358
rect 195980 245676 196032 245682
rect 195980 245618 196032 245624
rect 198004 245676 198056 245682
rect 198004 245618 198056 245624
rect 133604 243092 133656 243098
rect 133604 243034 133656 243040
rect 135904 243092 135956 243098
rect 135904 243034 135956 243040
rect 133616 242214 133644 243034
rect 124128 242208 124180 242214
rect 124128 242150 124180 242156
rect 133604 242208 133656 242214
rect 133604 242150 133656 242156
rect 124140 240854 124168 242150
rect 124128 240848 124180 240854
rect 124128 240790 124180 240796
rect 195992 240786 196020 245618
rect 195980 240780 196032 240786
rect 195980 240722 196032 240728
rect 50344 240576 50396 240582
rect 50344 240518 50396 240524
rect 395356 240106 395384 625806
rect 395344 240100 395396 240106
rect 395344 240042 395396 240048
rect 46848 239828 46900 239834
rect 46848 239770 46900 239776
rect 46756 239760 46808 239766
rect 46756 239702 46808 239708
rect 105820 233164 105872 233170
rect 105820 233106 105872 233112
rect 45744 232416 45796 232422
rect 45744 232358 45796 232364
rect 45836 232416 45888 232422
rect 45836 232358 45888 232364
rect 48320 232416 48372 232422
rect 48320 232358 48372 232364
rect 45756 231810 45784 232358
rect 46848 232348 46900 232354
rect 46848 232290 46900 232296
rect 45744 231804 45796 231810
rect 45744 231746 45796 231752
rect 46860 230450 46888 232290
rect 48332 230994 48360 232358
rect 105832 232014 105860 233106
rect 394700 232144 394752 232150
rect 394700 232086 394752 232092
rect 105820 232008 105872 232014
rect 105820 231950 105872 231956
rect 117964 232008 118016 232014
rect 117964 231950 118016 231956
rect 50620 231804 50672 231810
rect 50620 231746 50672 231752
rect 48320 230988 48372 230994
rect 48320 230930 48372 230936
rect 46940 230512 46992 230518
rect 46940 230454 46992 230460
rect 46848 230444 46900 230450
rect 46848 230386 46900 230392
rect 45652 230376 45704 230382
rect 45652 230318 45704 230324
rect 46952 225622 46980 230454
rect 49608 230444 49660 230450
rect 49608 230386 49660 230392
rect 49620 229094 49648 230386
rect 49620 229066 49740 229094
rect 49712 227526 49740 229066
rect 50632 227866 50660 231746
rect 72424 230988 72476 230994
rect 72424 230930 72476 230936
rect 51540 230376 51592 230382
rect 51540 230318 51592 230324
rect 50620 227860 50672 227866
rect 50620 227802 50672 227808
rect 49700 227520 49752 227526
rect 49700 227462 49752 227468
rect 46940 225616 46992 225622
rect 46940 225558 46992 225564
rect 51552 223650 51580 230318
rect 56508 227860 56560 227866
rect 56508 227802 56560 227808
rect 52368 227520 52420 227526
rect 52368 227462 52420 227468
rect 52380 224890 52408 227462
rect 56520 225282 56548 227802
rect 56508 225276 56560 225282
rect 56508 225218 56560 225224
rect 52380 224862 52500 224890
rect 51540 223644 51592 223650
rect 51540 223586 51592 223592
rect 52472 223514 52500 224862
rect 55864 223576 55916 223582
rect 55864 223518 55916 223524
rect 52460 223508 52512 223514
rect 52460 223450 52512 223456
rect 47584 220856 47636 220862
rect 47584 220798 47636 220804
rect 46204 216640 46256 216646
rect 46204 216582 46256 216588
rect 46216 209030 46244 216582
rect 47596 212498 47624 220798
rect 53840 217320 53892 217326
rect 53840 217262 53892 217268
rect 53852 214606 53880 217262
rect 53840 214600 53892 214606
rect 53840 214542 53892 214548
rect 55876 212498 55904 223518
rect 56048 223508 56100 223514
rect 56048 223450 56100 223456
rect 56060 220794 56088 223450
rect 56048 220788 56100 220794
rect 56048 220730 56100 220736
rect 47584 212492 47636 212498
rect 47584 212434 47636 212440
rect 52460 212492 52512 212498
rect 52460 212434 52512 212440
rect 55864 212492 55916 212498
rect 55864 212434 55916 212440
rect 46204 209024 46256 209030
rect 46204 208966 46256 208972
rect 48780 209024 48832 209030
rect 48780 208966 48832 208972
rect 48792 205630 48820 208966
rect 52472 208690 52500 212434
rect 52460 208684 52512 208690
rect 52460 208626 52512 208632
rect 55864 208684 55916 208690
rect 55864 208626 55916 208632
rect 48780 205624 48832 205630
rect 48780 205566 48832 205572
rect 55876 191826 55904 208626
rect 56416 205624 56468 205630
rect 56416 205566 56468 205572
rect 56428 202978 56456 205566
rect 56416 202972 56468 202978
rect 56416 202914 56468 202920
rect 56612 195974 56640 230588
rect 72436 227050 72464 230930
rect 72424 227044 72476 227050
rect 72424 226986 72476 226992
rect 77944 227044 77996 227050
rect 77944 226986 77996 226992
rect 57888 225616 57940 225622
rect 57888 225558 57940 225564
rect 57244 225276 57296 225282
rect 57244 225218 57296 225224
rect 57256 222222 57284 225218
rect 57900 222902 57928 225558
rect 57888 222896 57940 222902
rect 57888 222838 57940 222844
rect 65708 222896 65760 222902
rect 65708 222838 65760 222844
rect 57244 222216 57296 222222
rect 57244 222158 57296 222164
rect 60648 222148 60700 222154
rect 60648 222090 60700 222096
rect 56968 220788 57020 220794
rect 56968 220730 57020 220736
rect 56980 216510 57008 220730
rect 60660 219434 60688 222090
rect 65720 220794 65748 222838
rect 65708 220788 65760 220794
rect 65708 220730 65760 220736
rect 69388 220788 69440 220794
rect 69388 220730 69440 220736
rect 60660 219406 60780 219434
rect 56968 216504 57020 216510
rect 56968 216446 57020 216452
rect 59636 216504 59688 216510
rect 59636 216446 59688 216452
rect 59648 213246 59676 216446
rect 60752 213926 60780 219406
rect 69400 218074 69428 220730
rect 77956 218754 77984 226986
rect 77944 218748 77996 218754
rect 77944 218690 77996 218696
rect 69388 218068 69440 218074
rect 69388 218010 69440 218016
rect 71964 218000 72016 218006
rect 71964 217942 72016 217948
rect 71976 215354 72004 217942
rect 71964 215348 72016 215354
rect 71964 215290 72016 215296
rect 76564 215280 76616 215286
rect 76564 215222 76616 215228
rect 60740 213920 60792 213926
rect 60740 213862 60792 213868
rect 63500 213920 63552 213926
rect 63500 213862 63552 213868
rect 59636 213240 59688 213246
rect 59636 213182 59688 213188
rect 59268 212492 59320 212498
rect 59268 212434 59320 212440
rect 59280 209166 59308 212434
rect 63512 211070 63540 213862
rect 68284 213240 68336 213246
rect 68284 213182 68336 213188
rect 63500 211064 63552 211070
rect 63500 211006 63552 211012
rect 65892 211064 65944 211070
rect 65892 211006 65944 211012
rect 59268 209160 59320 209166
rect 59268 209102 59320 209108
rect 62120 209160 62172 209166
rect 62120 209102 62172 209108
rect 62132 205698 62160 209102
rect 65904 208418 65932 211006
rect 68296 208962 68324 213182
rect 68284 208956 68336 208962
rect 68284 208898 68336 208904
rect 75552 208956 75604 208962
rect 75552 208898 75604 208904
rect 65892 208412 65944 208418
rect 65892 208354 65944 208360
rect 71688 208344 71740 208350
rect 71688 208286 71740 208292
rect 71700 206938 71728 208286
rect 71700 206910 71820 206938
rect 62120 205692 62172 205698
rect 62120 205634 62172 205640
rect 66444 205624 66496 205630
rect 66444 205566 66496 205572
rect 62120 202972 62172 202978
rect 62120 202914 62172 202920
rect 62132 201482 62160 202914
rect 66456 201482 66484 205566
rect 71792 204270 71820 206910
rect 71780 204264 71832 204270
rect 71780 204206 71832 204212
rect 73804 204264 73856 204270
rect 73804 204206 73856 204212
rect 62120 201476 62172 201482
rect 62120 201418 62172 201424
rect 64236 201476 64288 201482
rect 64236 201418 64288 201424
rect 66444 201476 66496 201482
rect 66444 201418 66496 201424
rect 69664 201476 69716 201482
rect 69664 201418 69716 201424
rect 56600 195968 56652 195974
rect 56600 195910 56652 195916
rect 55864 191820 55916 191826
rect 55864 191762 55916 191768
rect 64144 191820 64196 191826
rect 64144 191762 64196 191768
rect 64156 171834 64184 191762
rect 64248 189786 64276 201418
rect 64236 189780 64288 189786
rect 64236 189722 64288 189728
rect 69676 186046 69704 201418
rect 73816 198286 73844 204206
rect 75564 201482 75592 208898
rect 76576 205426 76604 215222
rect 77944 214600 77996 214606
rect 77944 214542 77996 214548
rect 76564 205420 76616 205426
rect 76564 205362 76616 205368
rect 77956 201482 77984 214542
rect 78312 205420 78364 205426
rect 78312 205362 78364 205368
rect 75552 201476 75604 201482
rect 75552 201418 75604 201424
rect 76564 201476 76616 201482
rect 76564 201418 76616 201424
rect 77944 201476 77996 201482
rect 77944 201418 77996 201424
rect 73804 198280 73856 198286
rect 73804 198222 73856 198228
rect 75552 198280 75604 198286
rect 75552 198222 75604 198228
rect 75564 194682 75592 198222
rect 75552 194676 75604 194682
rect 75552 194618 75604 194624
rect 69756 189780 69808 189786
rect 69756 189722 69808 189728
rect 69664 186040 69716 186046
rect 69664 185982 69716 185988
rect 69768 175982 69796 189722
rect 76576 188222 76604 201418
rect 78324 201414 78352 205362
rect 80704 201476 80756 201482
rect 80704 201418 80756 201424
rect 78312 201408 78364 201414
rect 78312 201350 78364 201356
rect 79968 201408 80020 201414
rect 79968 201350 80020 201356
rect 79980 197402 80008 201350
rect 79968 197396 80020 197402
rect 79968 197338 80020 197344
rect 76656 194676 76708 194682
rect 76656 194618 76708 194624
rect 76564 188216 76616 188222
rect 76564 188158 76616 188164
rect 76668 187406 76696 194618
rect 78588 188216 78640 188222
rect 78588 188158 78640 188164
rect 76656 187400 76708 187406
rect 76656 187342 76708 187348
rect 78600 186266 78628 188158
rect 79968 187400 80020 187406
rect 79968 187342 80020 187348
rect 78600 186238 78720 186266
rect 71044 186040 71096 186046
rect 71044 185982 71096 185988
rect 71056 178362 71084 185982
rect 78692 184822 78720 186238
rect 79980 184890 80008 187342
rect 79968 184884 80020 184890
rect 79968 184826 80020 184832
rect 78680 184816 78732 184822
rect 78680 184758 78732 184764
rect 71044 178356 71096 178362
rect 71044 178298 71096 178304
rect 72424 178356 72476 178362
rect 72424 178298 72476 178304
rect 69756 175976 69808 175982
rect 69756 175918 69808 175924
rect 64144 171828 64196 171834
rect 64144 171770 64196 171776
rect 69940 171828 69992 171834
rect 69940 171770 69992 171776
rect 69952 168298 69980 171770
rect 69940 168292 69992 168298
rect 69940 168234 69992 168240
rect 72436 160478 72464 178298
rect 80716 168298 80744 201418
rect 84844 197328 84896 197334
rect 84844 197270 84896 197276
rect 84856 186998 84884 197270
rect 86972 195906 87000 230588
rect 115952 230574 116518 230602
rect 87512 218748 87564 218754
rect 87512 218690 87564 218696
rect 87524 209846 87552 218690
rect 87512 209840 87564 209846
rect 87512 209782 87564 209788
rect 95884 209840 95936 209846
rect 95884 209782 95936 209788
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 84844 186992 84896 186998
rect 84844 186934 84896 186940
rect 86224 186992 86276 186998
rect 86224 186934 86276 186940
rect 81440 184884 81492 184890
rect 81440 184826 81492 184832
rect 80796 184816 80848 184822
rect 80796 184758 80848 184764
rect 77208 168292 77260 168298
rect 77208 168234 77260 168240
rect 80704 168292 80756 168298
rect 80704 168234 80756 168240
rect 77220 164898 77248 168234
rect 80808 167074 80836 184758
rect 81452 182238 81480 184826
rect 81440 182232 81492 182238
rect 81440 182174 81492 182180
rect 86236 168910 86264 186934
rect 86316 182164 86368 182170
rect 86316 182106 86368 182112
rect 86328 173874 86356 182106
rect 92480 175976 92532 175982
rect 92480 175918 92532 175924
rect 86316 173868 86368 173874
rect 86316 173810 86368 173816
rect 87972 173868 88024 173874
rect 87972 173810 88024 173816
rect 87984 169862 88012 173810
rect 92492 171426 92520 175918
rect 92480 171420 92532 171426
rect 92480 171362 92532 171368
rect 94504 171420 94556 171426
rect 94504 171362 94556 171368
rect 87972 169856 88024 169862
rect 87972 169798 88024 169804
rect 88984 169856 89036 169862
rect 88984 169798 89036 169804
rect 86224 168904 86276 168910
rect 86224 168846 86276 168852
rect 88340 168904 88392 168910
rect 88340 168846 88392 168852
rect 86868 168292 86920 168298
rect 86868 168234 86920 168240
rect 80796 167068 80848 167074
rect 80796 167010 80848 167016
rect 82084 167068 82136 167074
rect 82084 167010 82136 167016
rect 77208 164892 77260 164898
rect 77208 164834 77260 164840
rect 72424 160472 72476 160478
rect 72424 160414 72476 160420
rect 76748 160472 76800 160478
rect 76748 160414 76800 160420
rect 76760 155922 76788 160414
rect 82096 158098 82124 167010
rect 85212 164892 85264 164898
rect 85212 164834 85264 164840
rect 85224 162858 85252 164834
rect 86880 164218 86908 168234
rect 88352 165578 88380 168846
rect 88340 165572 88392 165578
rect 88340 165514 88392 165520
rect 86868 164212 86920 164218
rect 86868 164154 86920 164160
rect 85212 162852 85264 162858
rect 85212 162794 85264 162800
rect 82084 158092 82136 158098
rect 82084 158034 82136 158040
rect 83464 158092 83516 158098
rect 83464 158034 83516 158040
rect 76748 155916 76800 155922
rect 76748 155858 76800 155864
rect 79324 155916 79376 155922
rect 79324 155858 79376 155864
rect 45560 147008 45612 147014
rect 45560 146950 45612 146956
rect 48964 147008 49016 147014
rect 48964 146950 49016 146956
rect 40040 141704 40092 141710
rect 40040 141646 40092 141652
rect 43444 139460 43496 139466
rect 43444 139402 43496 139408
rect 37924 121440 37976 121446
rect 37924 121382 37976 121388
rect 23480 117292 23532 117298
rect 23480 117234 23532 117240
rect 43456 111790 43484 139402
rect 48976 117978 49004 146950
rect 79336 140350 79364 155858
rect 79324 140344 79376 140350
rect 79324 140286 79376 140292
rect 82728 140344 82780 140350
rect 82728 140286 82780 140292
rect 82740 136626 82768 140286
rect 83476 140146 83504 158034
rect 88996 150482 89024 169798
rect 90364 165572 90416 165578
rect 90364 165514 90416 165520
rect 88984 150476 89036 150482
rect 88984 150418 89036 150424
rect 83464 140140 83516 140146
rect 83464 140082 83516 140088
rect 85028 140140 85080 140146
rect 85028 140082 85080 140088
rect 85040 138106 85068 140082
rect 90376 139874 90404 165514
rect 91560 164212 91612 164218
rect 91560 164154 91612 164160
rect 91572 159390 91600 164154
rect 91744 162852 91796 162858
rect 91744 162794 91796 162800
rect 91560 159384 91612 159390
rect 91560 159326 91612 159332
rect 91756 148374 91784 162794
rect 94516 160138 94544 171362
rect 94504 160132 94556 160138
rect 94504 160074 94556 160080
rect 94780 150408 94832 150414
rect 94780 150350 94832 150356
rect 91744 148368 91796 148374
rect 91744 148310 91796 148316
rect 94792 146334 94820 150350
rect 94780 146328 94832 146334
rect 94780 146270 94832 146276
rect 90364 139868 90416 139874
rect 90364 139810 90416 139816
rect 91468 139868 91520 139874
rect 91468 139810 91520 139816
rect 85028 138100 85080 138106
rect 85028 138042 85080 138048
rect 86224 138100 86276 138106
rect 86224 138042 86276 138048
rect 82740 136598 82860 136626
rect 82832 134910 82860 136598
rect 82820 134904 82872 134910
rect 82820 134846 82872 134852
rect 85212 134904 85264 134910
rect 85212 134846 85264 134852
rect 85224 126886 85252 134846
rect 86236 131170 86264 138042
rect 91480 135250 91508 139810
rect 91468 135244 91520 135250
rect 91468 135186 91520 135192
rect 93768 135244 93820 135250
rect 93768 135186 93820 135192
rect 93780 133770 93808 135186
rect 93780 133742 93900 133770
rect 86224 131164 86276 131170
rect 86224 131106 86276 131112
rect 89536 131164 89588 131170
rect 89536 131106 89588 131112
rect 89548 129674 89576 131106
rect 93872 130150 93900 133742
rect 93860 130144 93912 130150
rect 93860 130086 93912 130092
rect 95608 130144 95660 130150
rect 95608 130086 95660 130092
rect 89536 129668 89588 129674
rect 89536 129610 89588 129616
rect 92388 129668 92440 129674
rect 92388 129610 92440 129616
rect 85212 126880 85264 126886
rect 85212 126822 85264 126828
rect 88800 126880 88852 126886
rect 88800 126822 88852 126828
rect 88812 124098 88840 126822
rect 92400 125474 92428 129610
rect 95620 125526 95648 130086
rect 95608 125520 95660 125526
rect 92400 125446 92520 125474
rect 95608 125462 95660 125468
rect 88800 124092 88852 124098
rect 88800 124034 88852 124040
rect 92388 124092 92440 124098
rect 92388 124034 92440 124040
rect 92400 121786 92428 124034
rect 92492 123486 92520 125446
rect 92480 123480 92532 123486
rect 92480 123422 92532 123428
rect 92388 121780 92440 121786
rect 92388 121722 92440 121728
rect 94412 121780 94464 121786
rect 94412 121722 94464 121728
rect 94424 118318 94452 121722
rect 94412 118312 94464 118318
rect 94412 118254 94464 118260
rect 48964 117972 49016 117978
rect 48964 117914 49016 117920
rect 63500 117972 63552 117978
rect 63500 117914 63552 117920
rect 63512 114510 63540 117914
rect 95896 115938 95924 209782
rect 115952 194614 115980 230574
rect 117976 229770 118004 231950
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 179420 231192 179472 231198
rect 179420 231134 179472 231140
rect 159364 231056 159416 231062
rect 159364 230998 159416 231004
rect 146312 230574 146510 230602
rect 117964 229764 118016 229770
rect 117964 229706 118016 229712
rect 131764 229764 131816 229770
rect 131764 229706 131816 229712
rect 118792 228404 118844 228410
rect 118792 228346 118844 228352
rect 118700 218068 118752 218074
rect 118700 218010 118752 218016
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 115204 187740 115256 187746
rect 115204 187682 115256 187688
rect 98644 160064 98696 160070
rect 98644 160006 98696 160012
rect 98184 159384 98236 159390
rect 98184 159326 98236 159332
rect 98196 153202 98224 159326
rect 98184 153196 98236 153202
rect 98184 153138 98236 153144
rect 97264 146260 97316 146266
rect 97264 146202 97316 146208
rect 97276 128654 97304 146202
rect 98656 143546 98684 160006
rect 102784 153196 102836 153202
rect 102784 153138 102836 153144
rect 98644 143540 98696 143546
rect 98644 143482 98696 143488
rect 100944 143540 100996 143546
rect 100944 143482 100996 143488
rect 100956 140350 100984 143482
rect 102796 142866 102824 153138
rect 109684 148368 109736 148374
rect 109684 148310 109736 148316
rect 102784 142860 102836 142866
rect 102784 142802 102836 142808
rect 108304 142860 108356 142866
rect 108304 142802 108356 142808
rect 100944 140344 100996 140350
rect 100944 140286 100996 140292
rect 108316 133210 108344 142802
rect 108304 133204 108356 133210
rect 108304 133146 108356 133152
rect 97264 128648 97316 128654
rect 97264 128590 97316 128596
rect 99748 128648 99800 128654
rect 99748 128590 99800 128596
rect 97172 125520 97224 125526
rect 97172 125462 97224 125468
rect 97184 120902 97212 125462
rect 99760 124098 99788 128590
rect 109696 128382 109724 148310
rect 109684 128376 109736 128382
rect 109684 128318 109736 128324
rect 112444 128376 112496 128382
rect 112444 128318 112496 128324
rect 99748 124092 99800 124098
rect 99748 124034 99800 124040
rect 102048 124092 102100 124098
rect 102048 124034 102100 124040
rect 100760 123480 100812 123486
rect 100760 123422 100812 123428
rect 100772 121854 100800 123422
rect 100760 121848 100812 121854
rect 100760 121790 100812 121796
rect 97172 120896 97224 120902
rect 97172 120838 97224 120844
rect 102060 120018 102088 124034
rect 102140 121848 102192 121854
rect 102140 121790 102192 121796
rect 102048 120012 102100 120018
rect 102048 119954 102100 119960
rect 102152 118590 102180 121790
rect 105728 120896 105780 120902
rect 105728 120838 105780 120844
rect 104348 120012 104400 120018
rect 104348 119954 104400 119960
rect 102140 118584 102192 118590
rect 102140 118526 102192 118532
rect 104360 118454 104388 119954
rect 104716 118584 104768 118590
rect 104716 118526 104768 118532
rect 104348 118448 104400 118454
rect 104348 118390 104400 118396
rect 97172 118312 97224 118318
rect 97172 118254 97224 118260
rect 97184 116006 97212 118254
rect 97172 116000 97224 116006
rect 97172 115942 97224 115948
rect 95884 115932 95936 115938
rect 95884 115874 95936 115880
rect 98644 115932 98696 115938
rect 98644 115874 98696 115880
rect 100668 115932 100720 115938
rect 100668 115874 100720 115880
rect 63500 114504 63552 114510
rect 63500 114446 63552 114452
rect 43444 111784 43496 111790
rect 43444 111726 43496 111732
rect 98656 100706 98684 115874
rect 100680 111790 100708 115874
rect 104728 114442 104756 118526
rect 105740 115938 105768 120838
rect 112456 118590 112484 128318
rect 112444 118584 112496 118590
rect 112444 118526 112496 118532
rect 108304 118448 108356 118454
rect 108304 118390 108356 118396
rect 105728 115932 105780 115938
rect 105728 115874 105780 115880
rect 104716 114436 104768 114442
rect 104716 114378 104768 114384
rect 107936 114436 107988 114442
rect 107936 114378 107988 114384
rect 100668 111784 100720 111790
rect 100668 111726 100720 111732
rect 107948 110498 107976 114378
rect 107936 110492 107988 110498
rect 107936 110434 107988 110440
rect 98644 100700 98696 100706
rect 98644 100642 98696 100648
rect 100760 100700 100812 100706
rect 100760 100642 100812 100648
rect 100772 97306 100800 100642
rect 108316 98734 108344 118390
rect 110328 115932 110380 115938
rect 110328 115874 110380 115880
rect 110340 113150 110368 115874
rect 110328 113144 110380 113150
rect 110328 113086 110380 113092
rect 108304 98728 108356 98734
rect 108304 98670 108356 98676
rect 109684 98728 109736 98734
rect 109684 98670 109736 98676
rect 100760 97300 100812 97306
rect 100760 97242 100812 97248
rect 109696 93294 109724 98670
rect 109776 97300 109828 97306
rect 109776 97242 109828 97248
rect 109788 93634 109816 97242
rect 109776 93628 109828 93634
rect 109776 93570 109828 93576
rect 113824 93628 113876 93634
rect 113824 93570 113876 93576
rect 109684 93288 109736 93294
rect 109684 93230 109736 93236
rect 110420 93288 110472 93294
rect 110420 93230 110472 93236
rect 110432 91118 110460 93230
rect 110420 91112 110472 91118
rect 110420 91054 110472 91060
rect 113836 80714 113864 93570
rect 113824 80708 113876 80714
rect 113824 80650 113876 80656
rect 6918 79520 6974 79529
rect 115216 79490 115244 187682
rect 118332 144288 118384 144294
rect 118332 144230 118384 144236
rect 118240 144220 118292 144226
rect 118240 144162 118292 144168
rect 118148 141568 118200 141574
rect 118148 141510 118200 141516
rect 118056 140072 118108 140078
rect 118056 140014 118108 140020
rect 117318 136912 117374 136921
rect 117318 136847 117374 136856
rect 117332 136746 117360 136847
rect 117320 136740 117372 136746
rect 117320 136682 117372 136688
rect 117964 136196 118016 136202
rect 117964 136138 118016 136144
rect 117318 135416 117374 135425
rect 117318 135351 117374 135360
rect 117332 135318 117360 135351
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117320 133952 117372 133958
rect 117318 133920 117320 133929
rect 117372 133920 117374 133929
rect 117318 133855 117374 133864
rect 117780 133204 117832 133210
rect 117780 133146 117832 133152
rect 117320 132456 117372 132462
rect 117318 132424 117320 132433
rect 117372 132424 117374 132433
rect 117318 132359 117374 132368
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130937 117360 131038
rect 117318 130928 117374 130937
rect 117318 130863 117374 130872
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 129441 117360 129678
rect 117318 129432 117374 129441
rect 117318 129367 117374 129376
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127945 117360 128250
rect 117318 127936 117374 127945
rect 117318 127871 117374 127880
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 126449 117360 126890
rect 117318 126440 117374 126449
rect 117318 126375 117374 126384
rect 117320 125588 117372 125594
rect 117320 125530 117372 125536
rect 117332 124953 117360 125530
rect 117318 124944 117374 124953
rect 117318 124879 117374 124888
rect 117320 124160 117372 124166
rect 117320 124102 117372 124108
rect 117332 123457 117360 124102
rect 117318 123448 117374 123457
rect 117318 123383 117374 123392
rect 117792 122834 117820 133146
rect 117700 122806 117820 122834
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 121961 117360 122742
rect 117318 121952 117374 121961
rect 117318 121887 117374 121896
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 120465 117360 121382
rect 117318 120456 117374 120465
rect 117318 120391 117374 120400
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 118969 117360 120022
rect 117318 118960 117374 118969
rect 117318 118895 117374 118904
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 115480 118584 115532 118590
rect 115480 118526 115532 118532
rect 115492 115938 115520 118526
rect 117332 117473 117360 118594
rect 117318 117464 117374 117473
rect 117318 117399 117374 117408
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 115977 117360 117234
rect 117318 115968 117374 115977
rect 115480 115932 115532 115938
rect 117318 115903 117374 115912
rect 115480 115874 115532 115880
rect 117700 114510 117728 122806
rect 117976 118658 118004 136138
rect 117964 118652 118016 118658
rect 117964 118594 118016 118600
rect 118068 118538 118096 140014
rect 117884 118510 118096 118538
rect 117780 115932 117832 115938
rect 117780 115874 117832 115880
rect 117320 114504 117372 114510
rect 117318 114472 117320 114481
rect 117688 114504 117740 114510
rect 117372 114472 117374 114481
rect 117688 114446 117740 114452
rect 117318 114407 117374 114416
rect 117320 113144 117372 113150
rect 117320 113086 117372 113092
rect 117332 112985 117360 113086
rect 117318 112976 117374 112985
rect 117318 112911 117374 112920
rect 117320 111784 117372 111790
rect 117320 111726 117372 111732
rect 117332 111489 117360 111726
rect 117318 111480 117374 111489
rect 117318 111415 117374 111424
rect 117320 110424 117372 110430
rect 117320 110366 117372 110372
rect 117332 109993 117360 110366
rect 117318 109984 117374 109993
rect 117318 109919 117374 109928
rect 117792 97986 117820 115874
rect 117884 107001 117912 118510
rect 118056 118448 118108 118454
rect 118056 118390 118108 118396
rect 118068 108497 118096 118390
rect 118054 108488 118110 108497
rect 118054 108423 118110 108432
rect 117870 106992 117926 107001
rect 117870 106927 117926 106936
rect 118160 104009 118188 141510
rect 118146 104000 118202 104009
rect 118146 103935 118202 103944
rect 117780 97980 117832 97986
rect 117780 97922 117832 97928
rect 118252 95033 118280 144162
rect 118238 95024 118294 95033
rect 118238 94959 118294 94968
rect 118344 93537 118372 144230
rect 118516 142996 118568 143002
rect 118516 142938 118568 142944
rect 118424 142928 118476 142934
rect 118424 142870 118476 142876
rect 118330 93528 118386 93537
rect 118330 93463 118386 93472
rect 118436 92041 118464 142870
rect 118422 92032 118478 92041
rect 118422 91967 118478 91976
rect 115296 91044 115348 91050
rect 115296 90986 115348 90992
rect 6918 79455 6974 79464
rect 115204 79484 115256 79490
rect 115204 79426 115256 79432
rect 5080 78872 5132 78878
rect 5080 78814 5132 78820
rect 115308 78742 115336 90986
rect 118528 90545 118556 142938
rect 118608 139528 118660 139534
rect 118608 139470 118660 139476
rect 118514 90536 118570 90545
rect 118514 90471 118570 90480
rect 118620 86057 118648 139470
rect 118712 89049 118740 218010
rect 118804 101017 118832 228346
rect 131776 183462 131804 229706
rect 138664 227792 138716 227798
rect 138664 227734 138716 227740
rect 138676 196790 138704 227734
rect 146312 197418 146340 230574
rect 157984 228472 158036 228478
rect 157984 228414 158036 228420
rect 147772 202156 147824 202162
rect 147772 202098 147824 202104
rect 146142 197390 146340 197418
rect 147784 197404 147812 202098
rect 155960 199436 156012 199442
rect 155960 199378 156012 199384
rect 148968 198008 149020 198014
rect 148968 197950 149020 197956
rect 148980 197404 149008 197950
rect 155972 197470 156000 199378
rect 154488 197464 154540 197470
rect 154146 197412 154488 197418
rect 154146 197406 154540 197412
rect 155960 197464 156012 197470
rect 155960 197406 156012 197412
rect 154146 197390 154528 197406
rect 157996 197334 158024 228414
rect 159376 209846 159404 230998
rect 159364 209840 159416 209846
rect 159364 209782 159416 209788
rect 162124 209840 162176 209846
rect 162124 209782 162176 209788
rect 152740 197328 152792 197334
rect 152582 197276 152740 197282
rect 152582 197270 152792 197276
rect 157984 197328 158036 197334
rect 157984 197270 158036 197276
rect 152582 197254 152780 197270
rect 138664 196784 138716 196790
rect 138664 196726 138716 196732
rect 150926 196722 151216 196738
rect 150926 196716 151228 196722
rect 150926 196710 151176 196716
rect 151176 196658 151228 196664
rect 155960 196648 156012 196654
rect 155802 196596 155960 196602
rect 155802 196590 156012 196596
rect 155802 196574 156000 196590
rect 162136 196518 162164 209782
rect 176672 202162 176700 230588
rect 176660 202156 176712 202162
rect 176660 202098 176712 202104
rect 164240 196784 164292 196790
rect 164240 196726 164292 196732
rect 162124 196512 162176 196518
rect 162124 196454 162176 196460
rect 164148 196512 164200 196518
rect 164148 196454 164200 196460
rect 140424 196030 140530 196058
rect 157366 196030 157656 196058
rect 138112 195968 138164 195974
rect 138110 195936 138112 195945
rect 140424 195945 140452 196030
rect 138164 195936 138166 195945
rect 140410 195936 140466 195945
rect 138110 195871 138166 195880
rect 139400 195900 139452 195906
rect 157628 195906 157656 196030
rect 158824 195937 158852 196044
rect 160100 195968 160152 195974
rect 158810 195928 158866 195937
rect 140410 195871 140466 195880
rect 157616 195900 157668 195906
rect 139400 195842 139452 195848
rect 158810 195863 158866 195872
rect 160098 195936 160100 195945
rect 160152 195936 160154 195945
rect 160098 195871 160154 195880
rect 157616 195842 157668 195848
rect 139412 195537 139440 195842
rect 140778 195664 140834 195673
rect 140778 195599 140834 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 140792 194614 140820 195599
rect 140780 194608 140832 194614
rect 140780 194550 140832 194556
rect 164160 194546 164188 196454
rect 164148 194540 164200 194546
rect 164148 194482 164200 194488
rect 140870 191856 140926 191865
rect 140870 191791 140926 191800
rect 140778 191584 140834 191593
rect 140778 191519 140834 191528
rect 140792 184249 140820 191519
rect 140884 184385 140912 191791
rect 144366 191040 144422 191049
rect 144288 190998 144366 191026
rect 140962 190904 141018 190913
rect 140962 190839 141018 190848
rect 140870 184376 140926 184385
rect 140870 184311 140926 184320
rect 140778 184240 140834 184249
rect 140778 184175 140834 184184
rect 140976 184113 141004 190839
rect 140962 184104 141018 184113
rect 140962 184039 141018 184048
rect 131764 183456 131816 183462
rect 131764 183398 131816 183404
rect 133972 183456 134024 183462
rect 133972 183398 134024 183404
rect 121460 180192 121512 180198
rect 121460 180134 121512 180140
rect 118884 175976 118936 175982
rect 118884 175918 118936 175924
rect 118790 101008 118846 101017
rect 118790 100943 118846 100952
rect 118698 89040 118754 89049
rect 118698 88975 118754 88984
rect 118896 87553 118924 175918
rect 118976 164892 119028 164898
rect 118976 164834 119028 164840
rect 118988 98025 119016 164834
rect 119068 158024 119120 158030
rect 119068 157966 119120 157972
rect 118974 98016 119030 98025
rect 118974 97951 119030 97960
rect 119080 96529 119108 157966
rect 120724 142860 120776 142866
rect 120724 142802 120776 142808
rect 119252 141500 119304 141506
rect 119252 141442 119304 141448
rect 119160 141432 119212 141438
rect 119160 141374 119212 141380
rect 119172 99521 119200 141374
rect 119264 102513 119292 141442
rect 119988 140140 120040 140146
rect 119988 140082 120040 140088
rect 119344 136672 119396 136678
rect 119344 136614 119396 136620
rect 119250 102504 119306 102513
rect 119250 102439 119306 102448
rect 119158 99512 119214 99521
rect 119158 99447 119214 99456
rect 119066 96520 119122 96529
rect 119066 96455 119122 96464
rect 118882 87544 118938 87553
rect 118882 87479 118938 87488
rect 118606 86048 118662 86057
rect 118606 85983 118662 85992
rect 118514 83056 118570 83065
rect 118514 82991 118570 83000
rect 118422 81560 118478 81569
rect 118422 81495 118478 81504
rect 115296 78736 115348 78742
rect 115296 78678 115348 78684
rect 89720 78192 89772 78198
rect 89720 78134 89772 78140
rect 57244 78124 57296 78130
rect 57244 78066 57296 78072
rect 46204 78056 46256 78062
rect 46204 77998 46256 78004
rect 22744 77988 22796 77994
rect 22744 77930 22796 77936
rect 20718 76664 20774 76673
rect 20718 76599 20774 76608
rect 6920 75200 6972 75206
rect 6920 75142 6972 75148
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 16574 4200 18566
rect 6932 16574 6960 75142
rect 19340 42084 19392 42090
rect 19340 42026 19392 42032
rect 19352 16574 19380 42026
rect 20732 16574 20760 76599
rect 22098 43480 22154 43489
rect 22098 43415 22154 43424
rect 22112 16574 22140 43415
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4080 480 4108 4791
rect 5276 480 5304 16546
rect 6460 4956 6512 4962
rect 6460 4898 6512 4904
rect 6472 480 6500 4898
rect 7668 480 7696 16546
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 11152 10328 11204 10334
rect 11152 10270 11204 10276
rect 9956 7608 10008 7614
rect 9956 7550 10008 7556
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8772 480 8800 4762
rect 9968 480 9996 7550
rect 11164 480 11192 10270
rect 13544 4888 13596 4894
rect 13544 4830 13596 4836
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12360 480 12388 3946
rect 13556 480 13584 4830
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 15846
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15948 480 15976 5034
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 480 17080 3470
rect 18248 480 18276 6122
rect 19444 480 19472 16546
rect 20626 3360 20682 3369
rect 20626 3295 20682 3304
rect 20640 480 20668 3295
rect 21836 480 21864 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 4962 22784 77930
rect 44180 76628 44232 76634
rect 44180 76570 44232 76576
rect 30380 76560 30432 76566
rect 30380 76502 30432 76508
rect 27620 73908 27672 73914
rect 27620 73850 27672 73856
rect 26240 73840 26292 73846
rect 26240 73782 26292 73788
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 22744 4956 22796 4962
rect 22744 4898 22796 4904
rect 24216 4956 24268 4962
rect 24216 4898 24268 4904
rect 24228 480 24256 4898
rect 25332 480 25360 6258
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 73782
rect 27632 16574 27660 73850
rect 30392 16574 30420 76502
rect 35898 75304 35954 75313
rect 35898 75239 35954 75248
rect 42800 75268 42852 75274
rect 34520 44872 34572 44878
rect 34520 44814 34572 44820
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31772 16574 31800 18634
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27724 480 27752 16546
rect 28448 10396 28500 10402
rect 28448 10338 28500 10344
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 10338
rect 30104 1148 30156 1154
rect 30104 1090 30156 1096
rect 30116 480 30144 1090
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 33232 5024 33284 5030
rect 33232 4966 33284 4972
rect 33244 1154 33272 4966
rect 33232 1148 33284 1154
rect 33232 1090 33284 1096
rect 33612 480 33640 6190
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 44814
rect 35912 12434 35940 75239
rect 42800 75210 42852 75216
rect 40038 73808 40094 73817
rect 40038 73743 40094 73752
rect 40052 16574 40080 73743
rect 40052 16546 40264 16574
rect 39120 14476 39172 14482
rect 39120 14418 39172 14424
rect 35912 12406 36860 12434
rect 35992 10464 36044 10470
rect 35992 10406 36044 10412
rect 36004 480 36032 10406
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36832 354 36860 12406
rect 38382 7576 38438 7585
rect 38382 7511 38438 7520
rect 38396 480 38424 7511
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 14418
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41878 7712 41934 7721
rect 41878 7647 41934 7656
rect 41892 480 41920 7647
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 75210
rect 44192 16574 44220 76570
rect 45560 19984 45612 19990
rect 45560 19926 45612 19932
rect 45572 16574 45600 19926
rect 44192 16546 45048 16574
rect 45572 16546 46152 16574
rect 44272 7676 44324 7682
rect 44272 7618 44324 7624
rect 44284 480 44312 7618
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46124 3482 46152 16546
rect 46216 5098 46244 77998
rect 53838 75440 53894 75449
rect 51080 75404 51132 75410
rect 53838 75375 53894 75384
rect 51080 75346 51132 75352
rect 50160 9036 50212 9042
rect 50160 8978 50212 8984
rect 48964 7744 49016 7750
rect 48964 7686 49016 7692
rect 46204 5092 46256 5098
rect 46204 5034 46256 5040
rect 47860 3596 47912 3602
rect 47860 3538 47912 3544
rect 46124 3454 46704 3482
rect 46676 480 46704 3454
rect 47872 480 47900 3538
rect 48976 480 49004 7686
rect 50172 480 50200 8978
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 75346
rect 53852 16574 53880 75375
rect 53852 16546 54984 16574
rect 53748 9104 53800 9110
rect 53748 9046 53800 9052
rect 52552 5092 52604 5098
rect 52552 5034 52604 5040
rect 52564 480 52592 5034
rect 53760 480 53788 9046
rect 54956 480 54984 16546
rect 57150 8936 57206 8945
rect 57150 8871 57206 8880
rect 56046 7848 56102 7857
rect 56046 7783 56102 7792
rect 56060 480 56088 7783
rect 57164 3482 57192 8871
rect 57256 6322 57284 78066
rect 86960 76764 87012 76770
rect 86960 76706 87012 76712
rect 69020 76696 69072 76702
rect 69020 76638 69072 76644
rect 57978 75576 58034 75585
rect 57978 75511 58034 75520
rect 57992 16574 58020 75511
rect 64880 73976 64932 73982
rect 64880 73918 64932 73924
rect 64892 16574 64920 73918
rect 69032 16574 69060 76638
rect 78680 71052 78732 71058
rect 78680 70994 78732 71000
rect 70400 44940 70452 44946
rect 70400 44882 70452 44888
rect 70412 16574 70440 44882
rect 74540 22840 74592 22846
rect 74540 22782 74592 22788
rect 74552 16574 74580 22782
rect 78692 16574 78720 70994
rect 85580 20052 85632 20058
rect 85580 19994 85632 20000
rect 85592 16574 85620 19994
rect 86972 16574 87000 76706
rect 88340 36576 88392 36582
rect 88340 36518 88392 36524
rect 88352 16574 88380 36518
rect 89732 16574 89760 78134
rect 111798 76936 111854 76945
rect 111798 76871 111854 76880
rect 102140 76832 102192 76838
rect 93858 76800 93914 76809
rect 102140 76774 102192 76780
rect 93858 76735 93914 76744
rect 91098 44840 91154 44849
rect 91098 44775 91154 44784
rect 91112 16574 91140 44775
rect 57992 16546 58480 16574
rect 64892 16546 65104 16574
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 78692 16546 79272 16574
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 57244 6316 57296 6322
rect 57244 6258 57296 6264
rect 57164 3454 57284 3482
rect 57256 480 57284 3454
rect 58452 480 58480 16546
rect 64328 9308 64380 9314
rect 64328 9250 64380 9256
rect 63224 9240 63276 9246
rect 63224 9182 63276 9188
rect 60832 9172 60884 9178
rect 60832 9114 60884 9120
rect 59636 5160 59688 5166
rect 59636 5102 59688 5108
rect 59648 480 59676 5102
rect 60844 480 60872 9114
rect 62028 3664 62080 3670
rect 62028 3606 62080 3612
rect 62040 480 62068 3606
rect 63236 480 63264 9182
rect 64340 480 64368 9250
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 67916 9376 67968 9382
rect 67916 9318 67968 9324
rect 66720 6316 66772 6322
rect 66720 6258 66772 6264
rect 66732 480 66760 6258
rect 67928 480 67956 9318
rect 69112 3732 69164 3738
rect 69112 3674 69164 3680
rect 69124 480 69152 3674
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 73802 6216 73858 6225
rect 73802 6151 73858 6160
rect 72606 3496 72662 3505
rect 72606 3431 72662 3440
rect 72620 480 72648 3431
rect 73816 480 73844 6151
rect 75012 480 75040 16546
rect 78586 9072 78642 9081
rect 78586 9007 78642 9016
rect 77392 6384 77444 6390
rect 77392 6326 77444 6332
rect 76196 3800 76248 3806
rect 76196 3742 76248 3748
rect 76208 480 76236 3742
rect 77404 480 77432 6326
rect 78600 480 78628 9007
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 81624 10532 81676 10538
rect 81624 10474 81676 10480
rect 80888 6452 80940 6458
rect 80888 6394 80940 6400
rect 80900 480 80928 6394
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 10474
rect 84476 6520 84528 6526
rect 84476 6462 84528 6468
rect 83280 3868 83332 3874
rect 83280 3810 83332 3816
rect 83292 480 83320 3810
rect 84488 480 84516 6462
rect 85684 480 85712 16546
rect 86868 5228 86920 5234
rect 86868 5170 86920 5176
rect 86880 480 86908 5170
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92478 10296 92534 10305
rect 92478 10231 92534 10240
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10231
rect 93872 3466 93900 76735
rect 93952 74044 94004 74050
rect 93952 73986 94004 73992
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93964 480 93992 73986
rect 95240 53100 95292 53106
rect 95240 53042 95292 53048
rect 95252 16574 95280 53042
rect 95252 16546 95832 16574
rect 94780 3460 94832 3466
rect 94780 3402 94832 3408
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3402
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 99840 10600 99892 10606
rect 99840 10542 99892 10548
rect 98644 7812 98696 7818
rect 98644 7754 98696 7760
rect 97448 5296 97500 5302
rect 97448 5238 97500 5244
rect 97460 480 97488 5238
rect 98656 480 98684 7754
rect 99852 480 99880 10542
rect 102152 6914 102180 76774
rect 107660 75336 107712 75342
rect 107660 75278 107712 75284
rect 102232 65544 102284 65550
rect 102232 65486 102284 65492
rect 102244 16574 102272 65486
rect 107672 16574 107700 75278
rect 111812 16574 111840 76871
rect 118436 22778 118464 81495
rect 118528 60722 118556 82991
rect 119356 80034 119384 136614
rect 120000 136202 120028 140082
rect 119988 136196 120040 136202
rect 119988 136138 120040 136144
rect 120736 113174 120764 142802
rect 121276 140480 121328 140486
rect 121276 140422 121328 140428
rect 121288 138961 121316 140422
rect 121472 139890 121500 180134
rect 133984 180130 134012 183398
rect 136376 182022 136758 182050
rect 144288 182036 144316 190998
rect 144366 190975 144422 190984
rect 144460 190528 144512 190534
rect 144380 190476 144460 190482
rect 144380 190470 144512 190476
rect 144380 190454 144500 190470
rect 144380 182036 144408 190454
rect 145012 190324 145064 190330
rect 145012 190266 145064 190272
rect 145024 189106 145052 190266
rect 145852 189774 145958 189802
rect 144644 189100 144696 189106
rect 144644 189042 144696 189048
rect 145012 189100 145064 189106
rect 145012 189042 145064 189048
rect 136376 180198 136404 182022
rect 144656 181150 144684 189042
rect 145852 189009 145880 189774
rect 164252 189652 164280 196726
rect 167644 194540 167696 194546
rect 167644 194482 167696 194488
rect 145838 189000 145894 189009
rect 145838 188935 145894 188944
rect 144918 188184 144974 188193
rect 144918 188119 144974 188128
rect 144932 181257 144960 188119
rect 159560 185910 159588 188428
rect 159548 185904 159600 185910
rect 159548 185846 159600 185852
rect 159916 185564 159968 185570
rect 159916 185506 159968 185512
rect 144918 181248 144974 181257
rect 144918 181183 144974 181192
rect 144644 181144 144696 181150
rect 144644 181086 144696 181092
rect 151912 181076 151964 181082
rect 151912 181018 151964 181024
rect 144642 180976 144698 180985
rect 136468 180934 136758 180962
rect 144578 180934 144642 180962
rect 136364 180192 136416 180198
rect 136364 180134 136416 180140
rect 133972 180124 134024 180130
rect 133972 180066 134024 180072
rect 136468 178702 136496 180934
rect 144642 180911 144698 180920
rect 136560 179982 136758 180010
rect 122840 178696 122892 178702
rect 122840 178638 122892 178644
rect 136456 178696 136508 178702
rect 136456 178638 136508 178644
rect 122852 151814 122880 178638
rect 136364 178424 136416 178430
rect 136364 178366 136416 178372
rect 134984 177812 135036 177818
rect 134984 177754 135036 177760
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 124232 151814 124260 177278
rect 134996 176186 135024 177754
rect 135260 177268 135312 177274
rect 135260 177210 135312 177216
rect 126980 176180 127032 176186
rect 126980 176122 127032 176128
rect 134984 176180 135036 176186
rect 134984 176122 135036 176128
rect 125600 176044 125652 176050
rect 125600 175986 125652 175992
rect 125612 151814 125640 175986
rect 126992 151814 127020 176122
rect 135272 175234 135300 177210
rect 136376 176050 136404 178366
rect 136560 177970 136588 179982
rect 151924 179518 151952 181018
rect 159928 180742 159956 185506
rect 159916 180736 159968 180742
rect 159916 180678 159968 180684
rect 159916 180124 159968 180130
rect 159916 180066 159968 180072
rect 151912 179512 151964 179518
rect 151912 179454 151964 179460
rect 153936 179512 153988 179518
rect 157798 179480 157854 179489
rect 153988 179460 154436 179466
rect 153936 179454 154436 179460
rect 153948 179450 154436 179454
rect 149060 179444 149112 179450
rect 153948 179444 154448 179450
rect 153948 179438 154396 179444
rect 149060 179386 149112 179392
rect 157798 179415 157800 179424
rect 154396 179386 154448 179392
rect 157852 179415 157854 179424
rect 158534 179480 158590 179489
rect 158628 179444 158680 179450
rect 158590 179424 158628 179432
rect 158534 179415 158628 179424
rect 158548 179404 158628 179415
rect 157800 179386 157852 179392
rect 158628 179386 158680 179392
rect 136744 178838 136772 179044
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136732 178832 136784 178838
rect 136732 178774 136784 178780
rect 143078 178800 143134 178809
rect 143078 178735 143134 178744
rect 141606 178664 141662 178673
rect 141606 178599 141662 178608
rect 136468 177942 136588 177970
rect 136468 177342 136496 177942
rect 136744 177834 136772 177956
rect 136652 177818 136772 177834
rect 136640 177812 136772 177818
rect 136692 177806 136772 177812
rect 136640 177754 136692 177760
rect 136456 177336 136508 177342
rect 136456 177278 136508 177284
rect 136560 177274 136758 177290
rect 136548 177268 136758 177274
rect 136600 177262 136758 177268
rect 136548 177210 136600 177216
rect 136364 176044 136416 176050
rect 136364 175986 136416 175992
rect 136744 175794 136772 175916
rect 136560 175766 136772 175794
rect 128360 175228 128412 175234
rect 128360 175170 128412 175176
rect 135260 175228 135312 175234
rect 135260 175170 135312 175176
rect 128372 151814 128400 175170
rect 135904 174412 135956 174418
rect 135904 174354 135956 174360
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 131120 172576 131172 172582
rect 131120 172518 131172 172524
rect 122852 151786 122972 151814
rect 124232 151786 124536 151814
rect 125612 151786 126100 151814
rect 126992 151786 127664 151814
rect 128372 151786 129228 151814
rect 122840 143064 122892 143070
rect 122840 143006 122892 143012
rect 122852 140486 122880 143006
rect 122840 140480 122892 140486
rect 122840 140422 122892 140428
rect 122944 139890 122972 151786
rect 124508 139890 124536 151786
rect 126072 139890 126100 151786
rect 127636 139890 127664 151786
rect 129200 139890 129228 151786
rect 131132 139890 131160 172518
rect 132500 171148 132552 171154
rect 132500 171090 132552 171096
rect 132512 139890 132540 171090
rect 133892 139890 133920 173878
rect 135260 171692 135312 171698
rect 135260 171634 135312 171640
rect 135272 151814 135300 171634
rect 135272 151786 135484 151814
rect 134064 147688 134116 147694
rect 134064 147630 134116 147636
rect 134076 143070 134104 147630
rect 134064 143064 134116 143070
rect 134064 143006 134116 143012
rect 135456 139890 135484 151786
rect 135916 147694 135944 174354
rect 136560 172582 136588 175766
rect 136548 172576 136600 172582
rect 136548 172518 136600 172524
rect 136744 171154 136772 174964
rect 141620 174826 141648 178599
rect 141608 174820 141660 174826
rect 141608 174762 141660 174768
rect 143092 174758 143120 178735
rect 144104 176050 144132 178871
rect 144092 176044 144144 176050
rect 144092 175986 144144 175992
rect 144460 175840 144512 175846
rect 144460 175782 144512 175788
rect 143080 174752 143132 174758
rect 143080 174694 143132 174700
rect 137376 173936 137428 173942
rect 137428 173884 137586 173890
rect 137376 173878 137586 173884
rect 137388 173862 137586 173878
rect 138020 172168 138072 172174
rect 138020 172110 138072 172116
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 138032 151814 138060 172110
rect 138676 171698 138704 173196
rect 139596 173182 139702 173210
rect 138664 171692 138716 171698
rect 138664 171634 138716 171640
rect 138032 151786 138612 151814
rect 135904 147688 135956 147694
rect 135904 147630 135956 147636
rect 137744 143404 137796 143410
rect 137744 143346 137796 143352
rect 137756 139890 137784 143346
rect 121472 139862 121808 139890
rect 122944 139862 123372 139890
rect 124508 139862 124936 139890
rect 126072 139862 126500 139890
rect 127636 139862 128064 139890
rect 129200 139862 129628 139890
rect 131132 139862 131192 139890
rect 132512 139862 132756 139890
rect 133892 139862 134320 139890
rect 135456 139862 135884 139890
rect 137448 139862 137784 139890
rect 138584 139890 138612 151786
rect 139596 143410 139624 173182
rect 140792 172174 140820 173196
rect 140780 172168 140832 172174
rect 140780 172110 140832 172116
rect 141700 146260 141752 146266
rect 141700 146202 141752 146208
rect 139584 143404 139636 143410
rect 139584 143346 139636 143352
rect 140688 142180 140740 142186
rect 140688 142122 140740 142128
rect 140700 139890 140728 142122
rect 138584 139862 139012 139890
rect 140576 139862 140728 139890
rect 141712 139890 141740 146202
rect 142172 142186 142200 173196
rect 142632 161474 142660 173196
rect 143644 161474 143672 173196
rect 142448 161446 142660 161474
rect 143552 161446 143672 161474
rect 142448 146266 142476 161446
rect 142436 146260 142488 146266
rect 142436 146202 142488 146208
rect 142160 142180 142212 142186
rect 142160 142122 142212 142128
rect 143552 139890 143580 161446
rect 144472 143070 144500 175782
rect 149072 174826 149100 179386
rect 159928 176458 159956 180066
rect 159916 176452 159968 176458
rect 159916 176394 159968 176400
rect 149336 176044 149388 176050
rect 149336 175986 149388 175992
rect 149348 175681 149376 175986
rect 165068 175976 165120 175982
rect 163502 175944 163558 175953
rect 159180 175908 159232 175914
rect 165068 175918 165120 175924
rect 165158 175944 165214 175953
rect 163502 175879 163558 175888
rect 159180 175850 159232 175856
rect 149980 175840 150032 175846
rect 149980 175782 150032 175788
rect 149334 175672 149390 175681
rect 149334 175607 149390 175616
rect 149992 175508 150020 175782
rect 158168 175772 158220 175778
rect 158168 175714 158220 175720
rect 158180 175681 158208 175714
rect 158166 175672 158222 175681
rect 158166 175607 158222 175616
rect 159192 175438 159220 175850
rect 163516 175778 163544 175879
rect 165080 175817 165108 175918
rect 165158 175879 165160 175888
rect 165212 175879 165214 175888
rect 167000 175908 167052 175914
rect 165160 175850 165212 175856
rect 167000 175850 167052 175856
rect 163594 175808 163650 175817
rect 163504 175772 163556 175778
rect 163594 175743 163650 175752
rect 165066 175808 165122 175817
rect 165066 175743 165122 175752
rect 163504 175714 163556 175720
rect 163608 175710 163636 175743
rect 163596 175704 163648 175710
rect 163596 175646 163648 175652
rect 153936 175432 153988 175438
rect 154396 175432 154448 175438
rect 153988 175392 154396 175420
rect 153936 175374 153988 175380
rect 154396 175374 154448 175380
rect 159180 175432 159232 175438
rect 159180 175374 159232 175380
rect 155500 175296 155552 175302
rect 155500 175238 155552 175244
rect 146484 174820 146536 174826
rect 146484 174762 146536 174768
rect 149060 174820 149112 174826
rect 149060 174762 149112 174768
rect 146496 174350 146524 174762
rect 152372 174752 152424 174758
rect 152372 174694 152424 174700
rect 152384 174556 152412 174694
rect 155512 174554 155540 175238
rect 162492 174752 162544 174758
rect 162492 174694 162544 174700
rect 156512 174684 156564 174690
rect 156512 174626 156564 174632
rect 155500 174548 155552 174554
rect 155500 174490 155552 174496
rect 146484 174344 146536 174350
rect 146484 174286 146536 174292
rect 144460 143064 144512 143070
rect 144460 143006 144512 143012
rect 144932 139890 144960 173196
rect 146312 151814 146340 173196
rect 146680 161474 146708 173196
rect 146496 161446 146708 161474
rect 146312 151786 146432 151814
rect 146404 139890 146432 151786
rect 146496 143546 146524 161446
rect 146484 143540 146536 143546
rect 146484 143482 146536 143488
rect 147692 143478 147720 173196
rect 149348 172990 149376 173196
rect 149336 172984 149388 172990
rect 149336 172926 149388 172932
rect 149624 161474 149652 173196
rect 150440 172984 150492 172990
rect 150440 172926 150492 172932
rect 149532 161446 149652 161474
rect 148048 143540 148100 143546
rect 148048 143482 148100 143488
rect 147680 143472 147732 143478
rect 147680 143414 147732 143420
rect 148060 139890 148088 143482
rect 149532 142186 149560 161446
rect 149612 143472 149664 143478
rect 149612 143414 149664 143420
rect 149520 142180 149572 142186
rect 149520 142122 149572 142128
rect 149624 139890 149652 143414
rect 150452 142154 150480 172926
rect 150636 161474 150664 173196
rect 152660 161474 152688 173196
rect 150544 161446 150664 161474
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 150544 143138 150572 161446
rect 152476 143478 152504 161446
rect 153488 143546 153516 173182
rect 155222 171864 155278 171873
rect 155222 171799 155278 171808
rect 155236 164218 155264 171799
rect 155224 164212 155276 164218
rect 155224 164154 155276 164160
rect 153476 143540 153528 143546
rect 153476 143482 153528 143488
rect 152464 143472 152516 143478
rect 152464 143414 152516 143420
rect 150532 143132 150584 143138
rect 150532 143074 150584 143080
rect 154580 143132 154632 143138
rect 154580 143074 154632 143080
rect 152740 142180 152792 142186
rect 150452 142126 151124 142154
rect 151096 139890 151124 142126
rect 152740 142122 152792 142128
rect 152752 139890 152780 142122
rect 154592 139890 154620 143074
rect 156524 139890 156552 174626
rect 161480 174616 161532 174622
rect 161480 174558 161532 174564
rect 157352 142186 157380 173196
rect 160100 164212 160152 164218
rect 160100 164154 160152 164160
rect 160112 158098 160140 164154
rect 160100 158092 160152 158098
rect 160100 158034 160152 158040
rect 161492 151814 161520 174558
rect 162504 172938 162532 174694
rect 162504 172910 162900 172938
rect 162872 169998 162900 172910
rect 163516 170082 163544 175100
rect 163424 170054 163544 170082
rect 162860 169992 162912 169998
rect 162860 169934 162912 169940
rect 163424 161474 163452 170054
rect 163504 169992 163556 169998
rect 163504 169934 163556 169940
rect 163516 166274 163544 169934
rect 163608 166394 163636 173196
rect 164528 173182 164634 173210
rect 163596 166388 163648 166394
rect 163596 166330 163648 166336
rect 163516 166246 163728 166274
rect 163596 166184 163648 166190
rect 163596 166126 163648 166132
rect 163424 161446 163544 161474
rect 161492 151786 162072 151814
rect 158996 143540 159048 143546
rect 158996 143482 159048 143488
rect 157432 143472 157484 143478
rect 157432 143414 157484 143420
rect 157340 142180 157392 142186
rect 157340 142122 157392 142128
rect 141712 139862 142140 139890
rect 143552 139862 143704 139890
rect 144932 139862 145268 139890
rect 146404 139862 146832 139890
rect 148060 139862 148396 139890
rect 149624 139862 149960 139890
rect 151096 139862 151524 139890
rect 152752 139862 153088 139890
rect 154592 139862 154652 139890
rect 156216 139862 156552 139890
rect 157444 139890 157472 143414
rect 159008 139890 159036 143482
rect 160560 143064 160612 143070
rect 160560 143006 160612 143012
rect 160572 139890 160600 143006
rect 162044 139890 162072 151786
rect 163516 143070 163544 161446
rect 163608 143206 163636 166126
rect 163700 160138 163728 166246
rect 163688 160132 163740 160138
rect 163688 160074 163740 160080
rect 163596 143200 163648 143206
rect 163596 143142 163648 143148
rect 164528 143138 164556 173182
rect 165436 172984 165488 172990
rect 165436 172926 165488 172932
rect 164516 143132 164568 143138
rect 164516 143074 164568 143080
rect 163504 143064 163556 143070
rect 163504 143006 163556 143012
rect 163688 142180 163740 142186
rect 163688 142122 163740 142128
rect 163700 139890 163728 142122
rect 165448 139890 165476 172926
rect 166264 160132 166316 160138
rect 166264 160074 166316 160080
rect 166276 146946 166304 160074
rect 166356 158092 166408 158098
rect 166356 158034 166408 158040
rect 166368 147014 166396 158034
rect 166356 147008 166408 147014
rect 166356 146950 166408 146956
rect 166264 146940 166316 146946
rect 166264 146882 166316 146888
rect 167012 139890 167040 175850
rect 167656 173874 167684 194482
rect 169760 179444 169812 179450
rect 169760 179386 169812 179392
rect 167644 173868 167696 173874
rect 167644 173810 167696 173816
rect 169116 173868 169168 173874
rect 169116 173810 169168 173816
rect 169128 169794 169156 173810
rect 169116 169788 169168 169794
rect 169116 169730 169168 169736
rect 169772 151814 169800 179386
rect 170404 169788 170456 169794
rect 170404 169730 170456 169736
rect 170416 160750 170444 169730
rect 170404 160744 170456 160750
rect 170404 160686 170456 160692
rect 173900 160744 173952 160750
rect 173900 160686 173952 160692
rect 173912 157690 173940 160686
rect 173900 157684 173952 157690
rect 173900 157626 173952 157632
rect 175924 157684 175976 157690
rect 175924 157626 175976 157632
rect 169772 151786 169892 151814
rect 168380 147008 168432 147014
rect 168380 146950 168432 146956
rect 168392 139890 168420 146950
rect 169864 139890 169892 151786
rect 174636 143200 174688 143206
rect 174636 143142 174688 143148
rect 171506 142896 171562 142905
rect 171506 142831 171562 142840
rect 171520 139890 171548 142831
rect 173070 142760 173126 142769
rect 173070 142695 173126 142704
rect 173084 139890 173112 142695
rect 174648 139890 174676 143142
rect 175936 142186 175964 157626
rect 176200 143132 176252 143138
rect 176200 143074 176252 143080
rect 175924 142180 175976 142186
rect 175924 142122 175976 142128
rect 176212 139890 176240 143074
rect 178040 143064 178092 143070
rect 178040 143006 178092 143012
rect 178052 139890 178080 143006
rect 157444 139862 157780 139890
rect 159008 139862 159344 139890
rect 160572 139862 160908 139890
rect 162044 139862 162472 139890
rect 163700 139862 164036 139890
rect 165448 139862 165600 139890
rect 167012 139862 167164 139890
rect 168392 139862 168728 139890
rect 169864 139862 170292 139890
rect 171520 139862 171856 139890
rect 173084 139862 173420 139890
rect 174648 139862 174984 139890
rect 176212 139862 176548 139890
rect 178052 139862 178112 139890
rect 178224 139528 178276 139534
rect 178224 139470 178276 139476
rect 178236 139398 178264 139470
rect 178224 139392 178276 139398
rect 178224 139334 178276 139340
rect 121274 138952 121330 138961
rect 121274 138887 121330 138896
rect 179432 126177 179460 231134
rect 180800 231124 180852 231130
rect 180800 231066 180852 231072
rect 179512 213988 179564 213994
rect 179512 213930 179564 213936
rect 179524 132025 179552 213930
rect 180064 151836 180116 151842
rect 180064 151778 180116 151784
rect 179602 135552 179658 135561
rect 179602 135487 179658 135496
rect 179510 132016 179566 132025
rect 179510 131951 179566 131960
rect 179418 126168 179474 126177
rect 179418 126103 179474 126112
rect 120908 114504 120960 114510
rect 120908 114446 120960 114452
rect 120644 113146 120764 113174
rect 120644 106049 120672 113146
rect 120630 106040 120686 106049
rect 120630 105975 120686 105984
rect 120920 103514 120948 114446
rect 120736 103486 120948 103514
rect 120736 97730 120764 103486
rect 120920 97986 121040 98002
rect 120908 97980 121040 97986
rect 120960 97974 121040 97980
rect 120908 97922 120960 97928
rect 120736 97702 120948 97730
rect 120630 84280 120686 84289
rect 120448 84244 120500 84250
rect 120630 84215 120686 84224
rect 120448 84186 120500 84192
rect 119344 80028 119396 80034
rect 119344 79970 119396 79976
rect 120460 79150 120488 84186
rect 120644 81433 120672 84215
rect 120630 81424 120686 81433
rect 120630 81359 120686 81368
rect 120724 79620 120776 79626
rect 120724 79562 120776 79568
rect 120736 79422 120764 79562
rect 120724 79416 120776 79422
rect 120724 79358 120776 79364
rect 120448 79144 120500 79150
rect 120448 79086 120500 79092
rect 119988 78668 120040 78674
rect 119988 78610 120040 78616
rect 120000 76430 120028 78610
rect 120816 78328 120868 78334
rect 120816 78270 120868 78276
rect 119988 76424 120040 76430
rect 119988 76366 120040 76372
rect 120724 75812 120776 75818
rect 120724 75754 120776 75760
rect 118700 74112 118752 74118
rect 118700 74054 118752 74060
rect 118516 60716 118568 60722
rect 118516 60658 118568 60664
rect 118424 22772 118476 22778
rect 118424 22714 118476 22720
rect 117320 18760 117372 18766
rect 117320 18702 117372 18708
rect 102244 16546 103376 16574
rect 107672 16546 108160 16574
rect 111812 16546 112392 16574
rect 102152 6886 102272 6914
rect 101036 5364 101088 5370
rect 101036 5306 101088 5312
rect 101048 480 101076 5306
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 106464 10668 106516 10674
rect 106464 10610 106516 10616
rect 105728 7880 105780 7886
rect 105728 7822 105780 7828
rect 104532 6588 104584 6594
rect 104532 6530 104584 6536
rect 104544 480 104572 6530
rect 105740 480 105768 7822
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 10610
rect 108132 480 108160 16546
rect 110510 10432 110566 10441
rect 110510 10367 110566 10376
rect 109314 7984 109370 7993
rect 109314 7919 109370 7928
rect 109328 480 109356 7919
rect 110524 480 110552 10367
rect 111614 6352 111670 6361
rect 111614 6287 111670 6296
rect 111628 480 111656 6287
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 14544 114060 14550
rect 114008 14486 114060 14492
rect 114020 480 114048 14486
rect 116400 7948 116452 7954
rect 116400 7890 116452 7896
rect 115204 6656 115256 6662
rect 115204 6598 115256 6604
rect 115216 480 115244 6598
rect 116412 480 116440 7890
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117332 354 117360 18702
rect 118712 16574 118740 74054
rect 120080 40316 120132 40322
rect 120080 40258 120132 40264
rect 120092 16574 120120 40258
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 118804 480 118832 16546
rect 119896 4140 119948 4146
rect 119896 4082 119948 4088
rect 119908 480 119936 4082
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 14482 120764 75754
rect 120828 19990 120856 78270
rect 120920 77178 120948 97702
rect 120908 77172 120960 77178
rect 120908 77114 120960 77120
rect 121012 77110 121040 97974
rect 178960 82136 179012 82142
rect 178960 82078 179012 82084
rect 178406 81016 178462 81025
rect 178406 80951 178462 80960
rect 178314 80880 178370 80889
rect 178314 80815 178370 80824
rect 174728 80708 174780 80714
rect 174728 80650 174780 80656
rect 174544 80572 174596 80578
rect 174544 80514 174596 80520
rect 174452 80368 174504 80374
rect 174452 80310 174504 80316
rect 125048 80300 125100 80306
rect 125048 80242 125100 80248
rect 123668 80096 123720 80102
rect 123668 80038 123720 80044
rect 122932 79892 122984 79898
rect 122932 79834 122984 79840
rect 122944 77994 122972 79834
rect 123022 79792 123078 79801
rect 123022 79727 123078 79736
rect 122932 77988 122984 77994
rect 122932 77930 122984 77936
rect 122564 77716 122616 77722
rect 122564 77658 122616 77664
rect 121000 77104 121052 77110
rect 121000 77046 121052 77052
rect 122104 75880 122156 75886
rect 122104 75822 122156 75828
rect 121460 75472 121512 75478
rect 121460 75414 121512 75420
rect 120816 19984 120868 19990
rect 120816 19926 120868 19932
rect 121472 16574 121500 75414
rect 121472 16546 122052 16574
rect 120724 14476 120776 14482
rect 120724 14418 120776 14424
rect 122024 3482 122052 16546
rect 122116 4962 122144 75822
rect 122288 75676 122340 75682
rect 122288 75618 122340 75624
rect 122196 75540 122248 75546
rect 122196 75482 122248 75488
rect 122104 4956 122156 4962
rect 122104 4898 122156 4904
rect 122208 3670 122236 75482
rect 122300 18698 122328 75618
rect 122576 73846 122604 77658
rect 122840 76492 122892 76498
rect 122840 76434 122892 76440
rect 122564 73840 122616 73846
rect 122564 73782 122616 73788
rect 122288 18692 122340 18698
rect 122288 18634 122340 18640
rect 122852 16574 122880 76434
rect 123036 75206 123064 79727
rect 123484 77784 123536 77790
rect 123484 77726 123536 77732
rect 123024 75200 123076 75206
rect 123024 75142 123076 75148
rect 123496 40322 123524 77726
rect 123680 75313 123708 80038
rect 124956 79960 125008 79966
rect 124956 79902 125008 79908
rect 124864 76900 124916 76906
rect 124864 76842 124916 76848
rect 123666 75304 123722 75313
rect 123666 75239 123722 75248
rect 124772 74860 124824 74866
rect 124772 74802 124824 74808
rect 124784 70394 124812 74802
rect 124232 70366 124812 70394
rect 123484 40316 123536 40322
rect 123484 40258 123536 40264
rect 122852 16546 123064 16574
rect 122196 3664 122248 3670
rect 122196 3606 122248 3612
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124232 8974 124260 70366
rect 124312 21412 124364 21418
rect 124312 21354 124364 21360
rect 124324 16574 124352 21354
rect 124324 16546 124720 16574
rect 124220 8968 124272 8974
rect 124220 8910 124272 8916
rect 124692 480 124720 16546
rect 124876 4146 124904 76842
rect 124968 15910 124996 79902
rect 125060 36582 125088 80242
rect 174464 80238 174492 80310
rect 174556 80238 174584 80514
rect 174634 80336 174690 80345
rect 174634 80271 174636 80280
rect 174688 80271 174690 80280
rect 174636 80242 174688 80248
rect 174452 80232 174504 80238
rect 174452 80174 174504 80180
rect 174544 80232 174596 80238
rect 174544 80174 174596 80180
rect 125428 80022 125580 80050
rect 125324 79348 125376 79354
rect 125324 79290 125376 79296
rect 125336 78402 125364 79290
rect 125324 78396 125376 78402
rect 125324 78338 125376 78344
rect 125232 78260 125284 78266
rect 125232 78202 125284 78208
rect 125140 77988 125192 77994
rect 125140 77930 125192 77936
rect 125152 42090 125180 77930
rect 125244 53106 125272 78202
rect 125324 77920 125376 77926
rect 125324 77862 125376 77868
rect 125336 65550 125364 77862
rect 125428 74866 125456 80022
rect 125508 79824 125560 79830
rect 125508 79766 125560 79772
rect 125520 75954 125548 79766
rect 125658 79744 125686 80036
rect 125750 79937 125778 80036
rect 125736 79928 125792 79937
rect 125736 79863 125792 79872
rect 125658 79716 125732 79744
rect 125600 78396 125652 78402
rect 125600 78338 125652 78344
rect 125508 75948 125560 75954
rect 125508 75890 125560 75896
rect 125416 74860 125468 74866
rect 125416 74802 125468 74808
rect 125612 70394 125640 78338
rect 125704 76537 125732 79716
rect 125842 79676 125870 80036
rect 125934 79830 125962 80036
rect 126026 79898 126054 80036
rect 126118 79937 126146 80036
rect 126104 79928 126160 79937
rect 126014 79892 126066 79898
rect 126104 79863 126160 79872
rect 126014 79834 126066 79840
rect 125922 79824 125974 79830
rect 125922 79766 125974 79772
rect 126060 79756 126112 79762
rect 126210 79744 126238 80036
rect 126302 79898 126330 80036
rect 126394 79971 126422 80036
rect 126380 79962 126436 79971
rect 126290 79892 126342 79898
rect 126380 79897 126436 79906
rect 126290 79834 126342 79840
rect 126486 79778 126514 80036
rect 126578 79898 126606 80036
rect 126670 79898 126698 80036
rect 126762 79966 126790 80036
rect 126750 79960 126802 79966
rect 126750 79902 126802 79908
rect 126566 79892 126618 79898
rect 126566 79834 126618 79840
rect 126658 79892 126710 79898
rect 126658 79834 126710 79840
rect 126854 79812 126882 80036
rect 126946 79966 126974 80036
rect 127038 79966 127066 80036
rect 127130 79971 127158 80036
rect 126934 79960 126986 79966
rect 126934 79902 126986 79908
rect 127026 79960 127078 79966
rect 127026 79902 127078 79908
rect 127116 79962 127172 79971
rect 127116 79897 127172 79906
rect 126808 79784 126882 79812
rect 127072 79824 127124 79830
rect 126336 79756 126388 79762
rect 126210 79716 126284 79744
rect 126060 79698 126112 79704
rect 125796 79648 125870 79676
rect 125690 76528 125746 76537
rect 125690 76463 125746 76472
rect 125796 75993 125824 79648
rect 125876 79552 125928 79558
rect 125876 79494 125928 79500
rect 125968 79552 126020 79558
rect 125968 79494 126020 79500
rect 125782 75984 125838 75993
rect 125782 75919 125838 75928
rect 125612 70366 125824 70394
rect 125324 65544 125376 65550
rect 125324 65486 125376 65492
rect 125232 53100 125284 53106
rect 125232 53042 125284 53048
rect 125140 42084 125192 42090
rect 125140 42026 125192 42032
rect 125048 36576 125100 36582
rect 125048 36518 125100 36524
rect 124956 15904 125008 15910
rect 124956 15846 125008 15852
rect 125796 4826 125824 70366
rect 125888 4894 125916 79494
rect 125980 6186 126008 79494
rect 126072 7614 126100 79698
rect 126150 79656 126206 79665
rect 126150 79591 126206 79600
rect 126164 10334 126192 79591
rect 126256 79354 126284 79716
rect 126486 79750 126744 79778
rect 126336 79698 126388 79704
rect 126244 79348 126296 79354
rect 126244 79290 126296 79296
rect 126348 78062 126376 79698
rect 126336 78056 126388 78062
rect 126336 77998 126388 78004
rect 126336 77444 126388 77450
rect 126336 77386 126388 77392
rect 126244 75948 126296 75954
rect 126244 75890 126296 75896
rect 126256 18630 126284 75890
rect 126244 18624 126296 18630
rect 126244 18566 126296 18572
rect 126152 10328 126204 10334
rect 126152 10270 126204 10276
rect 126348 9314 126376 77386
rect 126428 72820 126480 72826
rect 126428 72762 126480 72768
rect 126336 9308 126388 9314
rect 126336 9250 126388 9256
rect 126060 7608 126112 7614
rect 126060 7550 126112 7556
rect 125968 6180 126020 6186
rect 125968 6122 126020 6128
rect 125876 4888 125928 4894
rect 125876 4830 125928 4836
rect 125784 4820 125836 4826
rect 125784 4762 125836 4768
rect 124864 4140 124916 4146
rect 124864 4082 124916 4088
rect 125876 4140 125928 4146
rect 125876 4082 125928 4088
rect 125888 480 125916 4082
rect 126440 3534 126468 72762
rect 126716 70394 126744 79750
rect 126808 72826 126836 79784
rect 127072 79766 127124 79772
rect 126980 79756 127032 79762
rect 126980 79698 127032 79704
rect 126888 79688 126940 79694
rect 126888 79630 126940 79636
rect 126900 73914 126928 79630
rect 126992 78130 127020 79698
rect 126980 78124 127032 78130
rect 126980 78066 127032 78072
rect 127084 77994 127112 79766
rect 127222 79676 127250 80036
rect 127314 79937 127342 80036
rect 127300 79928 127356 79937
rect 127300 79863 127356 79872
rect 127406 79744 127434 80036
rect 127498 79966 127526 80036
rect 127486 79960 127538 79966
rect 127486 79902 127538 79908
rect 127360 79716 127434 79744
rect 127590 79744 127618 80036
rect 127682 79898 127710 80036
rect 127774 79966 127802 80036
rect 127866 79971 127894 80036
rect 127762 79960 127814 79966
rect 127762 79902 127814 79908
rect 127852 79962 127908 79971
rect 127670 79892 127722 79898
rect 127852 79897 127908 79906
rect 127670 79834 127722 79840
rect 127714 79792 127770 79801
rect 127590 79716 127664 79744
rect 127958 79778 127986 80036
rect 128050 79966 128078 80036
rect 128142 79971 128170 80036
rect 128038 79960 128090 79966
rect 128038 79902 128090 79908
rect 128128 79962 128184 79971
rect 128234 79966 128262 80036
rect 128128 79897 128184 79906
rect 128222 79960 128274 79966
rect 128222 79902 128274 79908
rect 127714 79727 127770 79736
rect 127912 79750 127986 79778
rect 128084 79824 128136 79830
rect 128084 79766 128136 79772
rect 128176 79824 128228 79830
rect 128176 79766 128228 79772
rect 127222 79648 127296 79676
rect 127164 79552 127216 79558
rect 127164 79494 127216 79500
rect 127072 77988 127124 77994
rect 127072 77930 127124 77936
rect 126980 77852 127032 77858
rect 126980 77794 127032 77800
rect 126888 73908 126940 73914
rect 126888 73850 126940 73856
rect 126796 72820 126848 72826
rect 126796 72762 126848 72768
rect 126624 70366 126744 70394
rect 126624 4010 126652 70366
rect 126992 9042 127020 77794
rect 127070 44976 127126 44985
rect 127070 44911 127126 44920
rect 126980 9036 127032 9042
rect 126980 8978 127032 8984
rect 127084 6914 127112 44911
rect 127176 10402 127204 79494
rect 127268 76673 127296 79648
rect 127254 76664 127310 76673
rect 127254 76599 127310 76608
rect 127256 76288 127308 76294
rect 127256 76230 127308 76236
rect 127268 10470 127296 76230
rect 127360 75886 127388 79716
rect 127530 79656 127586 79665
rect 127530 79591 127586 79600
rect 127440 75948 127492 75954
rect 127440 75890 127492 75896
rect 127348 75880 127400 75886
rect 127348 75822 127400 75828
rect 127348 75744 127400 75750
rect 127348 75686 127400 75692
rect 127360 44878 127388 75686
rect 127348 44872 127400 44878
rect 127348 44814 127400 44820
rect 127256 10464 127308 10470
rect 127256 10406 127308 10412
rect 127164 10396 127216 10402
rect 127164 10338 127216 10344
rect 127084 6886 127388 6914
rect 126612 4004 126664 4010
rect 126612 3946 126664 3952
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 126428 3528 126480 3534
rect 126428 3470 126480 3476
rect 126992 480 127020 3538
rect 127360 3482 127388 6886
rect 127452 5030 127480 75890
rect 127544 6254 127572 79591
rect 127636 77722 127664 79716
rect 127624 77716 127676 77722
rect 127624 77658 127676 77664
rect 127624 76356 127676 76362
rect 127624 76298 127676 76304
rect 127532 6248 127584 6254
rect 127532 6190 127584 6196
rect 127440 5024 127492 5030
rect 127440 4966 127492 4972
rect 127636 3670 127664 76298
rect 127728 75954 127756 79727
rect 127912 76566 127940 79750
rect 127990 78160 128046 78169
rect 127990 78095 128046 78104
rect 127900 76560 127952 76566
rect 127900 76502 127952 76508
rect 127716 75948 127768 75954
rect 127716 75890 127768 75896
rect 128004 73817 128032 78095
rect 128096 75682 128124 79766
rect 128188 75750 128216 79766
rect 128326 79744 128354 80036
rect 128418 79966 128446 80036
rect 128510 79971 128538 80036
rect 128406 79960 128458 79966
rect 128406 79902 128458 79908
rect 128496 79962 128552 79971
rect 128496 79897 128552 79906
rect 128602 79778 128630 80036
rect 128694 79971 128722 80036
rect 128680 79962 128736 79971
rect 128680 79897 128736 79906
rect 128280 79716 128354 79744
rect 128556 79750 128630 79778
rect 128280 76294 128308 79716
rect 128556 79642 128584 79750
rect 128786 79744 128814 80036
rect 128878 79971 128906 80036
rect 128864 79962 128920 79971
rect 128864 79897 128920 79906
rect 128970 79898 128998 80036
rect 129062 79966 129090 80036
rect 129154 79966 129182 80036
rect 129050 79960 129102 79966
rect 129050 79902 129102 79908
rect 129142 79960 129194 79966
rect 129246 79937 129274 80036
rect 129338 79966 129366 80036
rect 129326 79960 129378 79966
rect 129142 79902 129194 79908
rect 129232 79928 129288 79937
rect 128958 79892 129010 79898
rect 129326 79902 129378 79908
rect 129430 79898 129458 80036
rect 129522 79898 129550 80036
rect 129614 79966 129642 80036
rect 129706 79966 129734 80036
rect 129798 79966 129826 80036
rect 129602 79960 129654 79966
rect 129602 79902 129654 79908
rect 129694 79960 129746 79966
rect 129694 79902 129746 79908
rect 129786 79960 129838 79966
rect 129786 79902 129838 79908
rect 129232 79863 129288 79872
rect 129418 79892 129470 79898
rect 128958 79834 129010 79840
rect 129418 79834 129470 79840
rect 129510 79892 129562 79898
rect 129510 79834 129562 79840
rect 129786 79824 129838 79830
rect 129706 79772 129786 79778
rect 129890 79812 129918 80036
rect 129982 79966 130010 80036
rect 129970 79960 130022 79966
rect 130074 79937 130102 80036
rect 129970 79902 130022 79908
rect 130060 79928 130116 79937
rect 130166 79898 130194 80036
rect 130258 79898 130286 80036
rect 130350 79937 130378 80036
rect 130336 79928 130392 79937
rect 130060 79863 130116 79872
rect 130154 79892 130206 79898
rect 130154 79834 130206 79840
rect 130246 79892 130298 79898
rect 130336 79863 130392 79872
rect 130246 79834 130298 79840
rect 129890 79784 130102 79812
rect 129706 79766 129838 79772
rect 130074 79778 130102 79784
rect 130442 79778 130470 80036
rect 130534 79966 130562 80036
rect 130522 79960 130574 79966
rect 130522 79902 130574 79908
rect 130626 79812 130654 80036
rect 128360 79620 128412 79626
rect 128360 79562 128412 79568
rect 128464 79614 128584 79642
rect 128740 79716 128814 79744
rect 128912 79756 128964 79762
rect 128372 76634 128400 79562
rect 128360 76628 128412 76634
rect 128360 76570 128412 76576
rect 128358 76528 128414 76537
rect 128358 76463 128414 76472
rect 128268 76288 128320 76294
rect 128268 76230 128320 76236
rect 128176 75744 128228 75750
rect 128176 75686 128228 75692
rect 128084 75676 128136 75682
rect 128084 75618 128136 75624
rect 128372 75274 128400 76463
rect 128464 75818 128492 79614
rect 128544 79552 128596 79558
rect 128544 79494 128596 79500
rect 128556 76702 128584 79494
rect 128636 78532 128688 78538
rect 128636 78474 128688 78480
rect 128544 76696 128596 76702
rect 128544 76638 128596 76644
rect 128452 75812 128504 75818
rect 128452 75754 128504 75760
rect 128648 75290 128676 78474
rect 128740 78033 128768 79716
rect 128912 79698 128964 79704
rect 129096 79756 129148 79762
rect 129096 79698 129148 79704
rect 129706 79750 129826 79766
rect 130074 79750 130148 79778
rect 128726 78024 128782 78033
rect 128726 77959 128782 77968
rect 128360 75268 128412 75274
rect 128360 75210 128412 75216
rect 128464 75262 128676 75290
rect 128728 75268 128780 75274
rect 128360 75064 128412 75070
rect 128360 75006 128412 75012
rect 127990 73808 128046 73817
rect 127990 73743 128046 73752
rect 128372 6914 128400 75006
rect 128464 22846 128492 75262
rect 128728 75210 128780 75216
rect 128544 75200 128596 75206
rect 128544 75142 128596 75148
rect 128452 22840 128504 22846
rect 128452 22782 128504 22788
rect 128556 7682 128584 75142
rect 128636 75132 128688 75138
rect 128636 75074 128688 75080
rect 128648 7750 128676 75074
rect 128740 9110 128768 75210
rect 128924 75206 128952 79698
rect 129108 78334 129136 79698
rect 129280 79688 129332 79694
rect 129186 79656 129242 79665
rect 129280 79630 129332 79636
rect 129372 79688 129424 79694
rect 129372 79630 129424 79636
rect 129706 79642 129734 79750
rect 129832 79688 129884 79694
rect 129186 79591 129242 79600
rect 129096 78328 129148 78334
rect 129096 78270 129148 78276
rect 129096 78056 129148 78062
rect 129096 77998 129148 78004
rect 129004 77988 129056 77994
rect 129004 77930 129056 77936
rect 128912 75200 128964 75206
rect 128912 75142 128964 75148
rect 128728 9104 128780 9110
rect 128728 9046 128780 9052
rect 128636 7744 128688 7750
rect 128636 7686 128688 7692
rect 128544 7676 128596 7682
rect 128544 7618 128596 7624
rect 128372 6886 128952 6914
rect 127624 3664 127676 3670
rect 127624 3606 127676 3612
rect 127360 3454 128216 3482
rect 128188 480 128216 3454
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 6886
rect 129016 3806 129044 77930
rect 129108 75410 129136 77998
rect 129200 76362 129228 79591
rect 129188 76356 129240 76362
rect 129188 76298 129240 76304
rect 129096 75404 129148 75410
rect 129096 75346 129148 75352
rect 129292 75138 129320 79630
rect 129384 77858 129412 79630
rect 129464 79620 129516 79626
rect 129464 79562 129516 79568
rect 129556 79620 129608 79626
rect 129706 79614 129780 79642
rect 129832 79630 129884 79636
rect 129924 79688 129976 79694
rect 129924 79630 129976 79636
rect 129556 79562 129608 79568
rect 129476 78062 129504 79562
rect 129464 78056 129516 78062
rect 129464 77998 129516 78004
rect 129372 77852 129424 77858
rect 129372 77794 129424 77800
rect 129372 77648 129424 77654
rect 129372 77590 129424 77596
rect 129280 75132 129332 75138
rect 129280 75074 129332 75080
rect 129384 70394 129412 77590
rect 129292 70366 129412 70394
rect 129568 70394 129596 79562
rect 129648 78056 129700 78062
rect 129752 78033 129780 79614
rect 129844 78062 129872 79630
rect 129832 78056 129884 78062
rect 129648 77998 129700 78004
rect 129738 78024 129794 78033
rect 129660 75274 129688 77998
rect 129832 77998 129884 78004
rect 129738 77959 129794 77968
rect 129740 77852 129792 77858
rect 129740 77794 129792 77800
rect 129648 75268 129700 75274
rect 129648 75210 129700 75216
rect 129752 73982 129780 77794
rect 129832 75744 129884 75750
rect 129832 75686 129884 75692
rect 129740 73976 129792 73982
rect 129740 73918 129792 73924
rect 129844 70394 129872 75686
rect 129568 70366 129688 70394
rect 129292 64874 129320 70366
rect 129108 64846 129320 64874
rect 129108 9178 129136 64846
rect 129096 9172 129148 9178
rect 129096 9114 129148 9120
rect 129660 5098 129688 70366
rect 129752 70366 129872 70394
rect 129752 16574 129780 70366
rect 129752 16546 129872 16574
rect 129648 5092 129700 5098
rect 129648 5034 129700 5040
rect 129004 3800 129056 3806
rect 129004 3742 129056 3748
rect 129844 3482 129872 16546
rect 129936 5166 129964 79630
rect 130016 79620 130068 79626
rect 130016 79562 130068 79568
rect 130028 78169 130056 79562
rect 130014 78160 130070 78169
rect 130014 78095 130070 78104
rect 130120 78033 130148 79750
rect 130200 79756 130252 79762
rect 130396 79750 130470 79778
rect 130580 79784 130654 79812
rect 130396 79744 130424 79750
rect 130200 79698 130252 79704
rect 130304 79716 130424 79744
rect 130106 78024 130162 78033
rect 130106 77959 130162 77968
rect 130212 77654 130240 79698
rect 130200 77648 130252 77654
rect 130200 77590 130252 77596
rect 130016 77512 130068 77518
rect 130016 77454 130068 77460
rect 130028 75750 130056 77454
rect 130304 75914 130332 79716
rect 130476 79688 130528 79694
rect 130396 79648 130476 79676
rect 130396 77450 130424 79648
rect 130476 79630 130528 79636
rect 130474 78024 130530 78033
rect 130474 77959 130530 77968
rect 130384 77444 130436 77450
rect 130384 77386 130436 77392
rect 130120 75886 130332 75914
rect 130016 75744 130068 75750
rect 130016 75686 130068 75692
rect 130016 75608 130068 75614
rect 130016 75550 130068 75556
rect 130028 6322 130056 75550
rect 130120 9246 130148 75886
rect 130488 75546 130516 77959
rect 130580 77858 130608 79784
rect 130718 79744 130746 80036
rect 130672 79716 130746 79744
rect 130568 77852 130620 77858
rect 130568 77794 130620 77800
rect 130672 75614 130700 79716
rect 130810 79676 130838 80036
rect 130902 79898 130930 80036
rect 130994 79966 131022 80036
rect 130982 79960 131034 79966
rect 130982 79902 131034 79908
rect 130890 79892 130942 79898
rect 130890 79834 130942 79840
rect 130936 79756 130988 79762
rect 131086 79744 131114 80036
rect 131178 79898 131206 80036
rect 131270 79971 131298 80036
rect 131256 79962 131312 79971
rect 131166 79892 131218 79898
rect 131256 79897 131312 79906
rect 131362 79898 131390 80036
rect 131454 79971 131482 80036
rect 131440 79962 131496 79971
rect 131546 79966 131574 80036
rect 131638 79971 131666 80036
rect 131166 79834 131218 79840
rect 131350 79892 131402 79898
rect 131440 79897 131496 79906
rect 131534 79960 131586 79966
rect 131534 79902 131586 79908
rect 131624 79962 131680 79971
rect 131730 79966 131758 80036
rect 131624 79897 131680 79906
rect 131718 79960 131770 79966
rect 131718 79902 131770 79908
rect 131350 79834 131402 79840
rect 131822 79830 131850 80036
rect 131914 79971 131942 80036
rect 131900 79962 131956 79971
rect 131900 79897 131956 79906
rect 132006 79898 132034 80036
rect 131994 79892 132046 79898
rect 131994 79834 132046 79840
rect 131488 79824 131540 79830
rect 131394 79792 131450 79801
rect 131086 79716 131160 79744
rect 131488 79766 131540 79772
rect 131810 79824 131862 79830
rect 131810 79766 131862 79772
rect 131394 79727 131450 79736
rect 130936 79698 130988 79704
rect 130764 79648 130838 79676
rect 130660 75608 130712 75614
rect 130660 75550 130712 75556
rect 130476 75540 130528 75546
rect 130476 75482 130528 75488
rect 130764 75426 130792 79648
rect 130948 75914 130976 79698
rect 131028 79552 131080 79558
rect 131028 79494 131080 79500
rect 131040 78033 131068 79494
rect 131026 78024 131082 78033
rect 131026 77959 131082 77968
rect 131132 75914 131160 79716
rect 131212 79688 131264 79694
rect 131212 79630 131264 79636
rect 131224 78538 131252 79630
rect 131212 78532 131264 78538
rect 131212 78474 131264 78480
rect 131212 78328 131264 78334
rect 131212 78270 131264 78276
rect 130212 75398 130792 75426
rect 130856 75886 130976 75914
rect 131040 75886 131160 75914
rect 131224 75914 131252 78270
rect 131408 77994 131436 79727
rect 131396 77988 131448 77994
rect 131396 77930 131448 77936
rect 131224 75886 131344 75914
rect 130212 9382 130240 75398
rect 130292 75268 130344 75274
rect 130292 75210 130344 75216
rect 130304 44946 130332 75210
rect 130382 74488 130438 74497
rect 130382 74423 130438 74432
rect 130292 44940 130344 44946
rect 130292 44882 130344 44888
rect 130200 9376 130252 9382
rect 130200 9318 130252 9324
rect 130108 9240 130160 9246
rect 130108 9182 130160 9188
rect 130016 6316 130068 6322
rect 130016 6258 130068 6264
rect 129924 5160 129976 5166
rect 129924 5102 129976 5108
rect 130396 3602 130424 74423
rect 130856 70394 130884 75886
rect 131040 75274 131068 75886
rect 131028 75268 131080 75274
rect 131028 75210 131080 75216
rect 130764 70366 130884 70394
rect 130764 64874 130792 70366
rect 130580 64846 130792 64874
rect 130580 16574 130608 64846
rect 130580 16546 130700 16574
rect 130672 3738 130700 16546
rect 131316 6526 131344 75886
rect 131500 75290 131528 79766
rect 131672 79756 131724 79762
rect 132098 79744 132126 80036
rect 131672 79698 131724 79704
rect 131960 79716 132126 79744
rect 131580 78736 131632 78742
rect 131580 78678 131632 78684
rect 131592 75342 131620 78678
rect 131684 77586 131712 79698
rect 131764 79688 131816 79694
rect 131764 79630 131816 79636
rect 131854 79656 131910 79665
rect 131672 77580 131724 77586
rect 131672 77522 131724 77528
rect 131408 75262 131528 75290
rect 131580 75336 131632 75342
rect 131580 75278 131632 75284
rect 131304 6520 131356 6526
rect 131304 6462 131356 6468
rect 131408 6390 131436 75262
rect 131776 75154 131804 79630
rect 131854 79591 131910 79600
rect 131500 75126 131804 75154
rect 131500 6458 131528 75126
rect 131868 75018 131896 79591
rect 131960 78334 131988 79716
rect 132040 79552 132092 79558
rect 132190 79540 132218 80036
rect 132282 79898 132310 80036
rect 132374 79971 132402 80036
rect 132360 79962 132416 79971
rect 132270 79892 132322 79898
rect 132360 79897 132416 79906
rect 132466 79898 132494 80036
rect 132270 79834 132322 79840
rect 132454 79892 132506 79898
rect 132454 79834 132506 79840
rect 132558 79830 132586 80036
rect 132650 79971 132678 80036
rect 132636 79962 132692 79971
rect 132636 79897 132692 79906
rect 132546 79824 132598 79830
rect 132314 79792 132370 79801
rect 132546 79766 132598 79772
rect 132314 79727 132370 79736
rect 132742 79744 132770 80036
rect 132834 79898 132862 80036
rect 132926 79966 132954 80036
rect 132914 79960 132966 79966
rect 132914 79902 132966 79908
rect 132822 79892 132874 79898
rect 132822 79834 132874 79840
rect 132040 79494 132092 79500
rect 132144 79512 132218 79540
rect 131948 78328 132000 78334
rect 131948 78270 132000 78276
rect 132052 78112 132080 79494
rect 131592 74990 131896 75018
rect 131960 78084 132080 78112
rect 131592 10538 131620 74990
rect 131672 74928 131724 74934
rect 131672 74870 131724 74876
rect 131684 20058 131712 74870
rect 131960 70394 131988 78084
rect 132040 77580 132092 77586
rect 132040 77522 132092 77528
rect 132052 71058 132080 77522
rect 132144 74934 132172 79512
rect 132224 77988 132276 77994
rect 132224 77930 132276 77936
rect 132132 74928 132184 74934
rect 132132 74870 132184 74876
rect 132040 71052 132092 71058
rect 132040 70994 132092 71000
rect 132236 70394 132264 77930
rect 132328 76770 132356 79727
rect 132742 79716 132816 79744
rect 132408 79688 132460 79694
rect 132788 79676 132816 79716
rect 133018 79676 133046 80036
rect 133110 79744 133138 80036
rect 133202 79898 133230 80036
rect 133190 79892 133242 79898
rect 133190 79834 133242 79840
rect 133110 79716 133184 79744
rect 132408 79630 132460 79636
rect 132498 79656 132554 79665
rect 132420 78198 132448 79630
rect 132788 79648 132908 79676
rect 132498 79591 132554 79600
rect 132592 79620 132644 79626
rect 132408 78192 132460 78198
rect 132408 78134 132460 78140
rect 132512 76838 132540 79591
rect 132592 79562 132644 79568
rect 132500 76832 132552 76838
rect 132604 76809 132632 79562
rect 132684 79552 132736 79558
rect 132684 79494 132736 79500
rect 132776 79552 132828 79558
rect 132776 79494 132828 79500
rect 132696 77994 132724 79494
rect 132684 77988 132736 77994
rect 132684 77930 132736 77936
rect 132788 77722 132816 79494
rect 132776 77716 132828 77722
rect 132776 77658 132828 77664
rect 132880 77489 132908 79648
rect 132972 79648 133046 79676
rect 132972 78266 133000 79648
rect 133052 79552 133104 79558
rect 133052 79494 133104 79500
rect 132960 78260 133012 78266
rect 132960 78202 133012 78208
rect 133064 77976 133092 79494
rect 132972 77948 133092 77976
rect 132866 77480 132922 77489
rect 132866 77415 132922 77424
rect 132500 76774 132552 76780
rect 132590 76800 132646 76809
rect 132316 76764 132368 76770
rect 132590 76735 132646 76744
rect 132316 76706 132368 76712
rect 132592 76696 132644 76702
rect 132592 76638 132644 76644
rect 131868 70366 131988 70394
rect 132052 70366 132264 70394
rect 131672 20052 131724 20058
rect 131672 19994 131724 20000
rect 131580 10532 131632 10538
rect 131580 10474 131632 10480
rect 131488 6452 131540 6458
rect 131488 6394 131540 6400
rect 131396 6384 131448 6390
rect 131396 6326 131448 6332
rect 131868 3874 131896 70366
rect 132052 5234 132080 70366
rect 132604 5302 132632 76638
rect 132972 75914 133000 77948
rect 133052 77852 133104 77858
rect 133052 77794 133104 77800
rect 132788 75886 133000 75914
rect 132684 75336 132736 75342
rect 132684 75278 132736 75284
rect 132696 6594 132724 75278
rect 132788 7818 132816 75886
rect 132868 75268 132920 75274
rect 132868 75210 132920 75216
rect 132880 7886 132908 75210
rect 132960 75200 133012 75206
rect 132960 75142 133012 75148
rect 132972 10674 133000 75142
rect 132960 10668 133012 10674
rect 132960 10610 133012 10616
rect 133064 10606 133092 77794
rect 133156 76702 133184 79716
rect 133294 79676 133322 80036
rect 133386 79830 133414 80036
rect 133478 79903 133506 80036
rect 133464 79894 133520 79903
rect 133374 79824 133426 79830
rect 133464 79829 133520 79838
rect 133570 79778 133598 80036
rect 133662 79830 133690 80036
rect 133754 79898 133782 80036
rect 133846 79937 133874 80036
rect 133938 79966 133966 80036
rect 133926 79960 133978 79966
rect 133832 79928 133888 79937
rect 133742 79892 133794 79898
rect 133926 79902 133978 79908
rect 133832 79863 133888 79872
rect 133742 79834 133794 79840
rect 133374 79766 133426 79772
rect 133478 79750 133598 79778
rect 133650 79824 133702 79830
rect 133650 79766 133702 79772
rect 133880 79824 133932 79830
rect 134030 79801 134058 80036
rect 134122 79966 134150 80036
rect 134214 79971 134242 80036
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 134200 79962 134256 79971
rect 134306 79966 134334 80036
rect 134398 79971 134426 80036
rect 134200 79897 134256 79906
rect 134294 79960 134346 79966
rect 134294 79902 134346 79908
rect 134384 79962 134440 79971
rect 134384 79897 134440 79906
rect 133880 79766 133932 79772
rect 134016 79792 134072 79801
rect 133478 79676 133506 79750
rect 133248 79648 133322 79676
rect 133432 79648 133506 79676
rect 133786 79656 133842 79665
rect 133248 77858 133276 79648
rect 133328 79552 133380 79558
rect 133328 79494 133380 79500
rect 133236 77852 133288 77858
rect 133236 77794 133288 77800
rect 133236 77716 133288 77722
rect 133236 77658 133288 77664
rect 133144 76696 133196 76702
rect 133144 76638 133196 76644
rect 133248 74050 133276 77658
rect 133236 74044 133288 74050
rect 133236 73986 133288 73992
rect 133340 70394 133368 79494
rect 133432 77926 133460 79648
rect 133604 79620 133656 79626
rect 133786 79591 133842 79600
rect 133604 79562 133656 79568
rect 133420 77920 133472 77926
rect 133420 77862 133472 77868
rect 133512 77444 133564 77450
rect 133512 77386 133564 77392
rect 133156 70366 133368 70394
rect 133524 70394 133552 77386
rect 133616 75342 133644 79562
rect 133696 79552 133748 79558
rect 133696 79494 133748 79500
rect 133604 75336 133656 75342
rect 133604 75278 133656 75284
rect 133708 75274 133736 79494
rect 133696 75268 133748 75274
rect 133696 75210 133748 75216
rect 133800 75206 133828 79591
rect 133892 78742 133920 79766
rect 134016 79727 134072 79736
rect 134338 79792 134394 79801
rect 134338 79727 134394 79736
rect 134490 79744 134518 80036
rect 134582 79898 134610 80036
rect 134570 79892 134622 79898
rect 134570 79834 134622 79840
rect 134674 79744 134702 80036
rect 134766 79898 134794 80036
rect 134858 79937 134886 80036
rect 134844 79928 134900 79937
rect 134754 79892 134806 79898
rect 134844 79863 134900 79872
rect 134754 79834 134806 79840
rect 134798 79792 134854 79801
rect 134064 79688 134116 79694
rect 134062 79656 134064 79665
rect 134116 79656 134118 79665
rect 134062 79591 134118 79600
rect 134156 79620 134208 79626
rect 134156 79562 134208 79568
rect 133972 79552 134024 79558
rect 133972 79494 134024 79500
rect 133880 78736 133932 78742
rect 133880 78678 133932 78684
rect 133984 78282 134012 79494
rect 134064 79484 134116 79490
rect 134064 79426 134116 79432
rect 134076 78878 134104 79426
rect 134064 78872 134116 78878
rect 134064 78814 134116 78820
rect 133984 78254 134104 78282
rect 133972 78192 134024 78198
rect 133972 78134 134024 78140
rect 133880 77988 133932 77994
rect 133880 77930 133932 77936
rect 133788 75200 133840 75206
rect 133788 75142 133840 75148
rect 133524 70366 133828 70394
rect 133052 10600 133104 10606
rect 133052 10542 133104 10548
rect 132868 7880 132920 7886
rect 132868 7822 132920 7828
rect 132776 7812 132828 7818
rect 132776 7754 132828 7760
rect 132684 6588 132736 6594
rect 132684 6530 132736 6536
rect 133156 5370 133184 70366
rect 133144 5364 133196 5370
rect 133144 5306 133196 5312
rect 132592 5296 132644 5302
rect 132592 5238 132644 5244
rect 132040 5228 132092 5234
rect 132040 5170 132092 5176
rect 131856 3868 131908 3874
rect 131856 3810 131908 3816
rect 131764 3800 131816 3806
rect 131764 3742 131816 3748
rect 130660 3732 130712 3738
rect 130660 3674 130712 3680
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 129844 3454 130608 3482
rect 130580 480 130608 3454
rect 131776 480 131804 3742
rect 132960 3664 133012 3670
rect 132960 3606 133012 3612
rect 132972 480 133000 3606
rect 133800 3534 133828 70366
rect 133788 3528 133840 3534
rect 133788 3470 133840 3476
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 77930
rect 133984 70394 134012 78134
rect 134076 74118 134104 78254
rect 134168 76945 134196 79562
rect 134154 76936 134210 76945
rect 134154 76871 134210 76880
rect 134352 75914 134380 79727
rect 134490 79716 134564 79744
rect 134674 79716 134748 79744
rect 134950 79744 134978 80036
rect 135042 79966 135070 80036
rect 135134 79966 135162 80036
rect 135030 79960 135082 79966
rect 135030 79902 135082 79908
rect 135122 79960 135174 79966
rect 135122 79902 135174 79908
rect 135226 79812 135254 80036
rect 135318 79830 135346 80036
rect 135410 79937 135438 80036
rect 135502 79966 135530 80036
rect 135490 79960 135542 79966
rect 135396 79928 135452 79937
rect 135490 79902 135542 79908
rect 135396 79863 135452 79872
rect 134798 79727 134854 79736
rect 134432 79620 134484 79626
rect 134432 79562 134484 79568
rect 134444 78198 134472 79562
rect 134536 79472 134564 79716
rect 134536 79444 134656 79472
rect 134524 79348 134576 79354
rect 134524 79290 134576 79296
rect 134432 78192 134484 78198
rect 134432 78134 134484 78140
rect 134432 78056 134484 78062
rect 134432 77998 134484 78004
rect 134168 75886 134380 75914
rect 134064 74112 134116 74118
rect 134064 74054 134116 74060
rect 133984 70366 134104 70394
rect 134076 7954 134104 70366
rect 134168 14550 134196 75886
rect 134248 75268 134300 75274
rect 134248 75210 134300 75216
rect 134260 18766 134288 75210
rect 134444 70394 134472 77998
rect 134352 70366 134472 70394
rect 134352 21418 134380 70366
rect 134340 21412 134392 21418
rect 134340 21354 134392 21360
rect 134248 18760 134300 18766
rect 134248 18702 134300 18708
rect 134156 14544 134208 14550
rect 134156 14486 134208 14492
rect 134064 7948 134116 7954
rect 134064 7890 134116 7896
rect 134536 4146 134564 79290
rect 134628 70394 134656 79444
rect 134720 75274 134748 79716
rect 134812 76906 134840 79727
rect 134904 79716 134978 79744
rect 135180 79784 135254 79812
rect 135306 79824 135358 79830
rect 134904 77790 134932 79716
rect 134984 79620 135036 79626
rect 134984 79562 135036 79568
rect 135076 79620 135128 79626
rect 135076 79562 135128 79568
rect 134892 77784 134944 77790
rect 134892 77726 134944 77732
rect 134800 76900 134852 76906
rect 134800 76842 134852 76848
rect 134996 75478 135024 79562
rect 135088 76498 135116 79562
rect 135180 78062 135208 79784
rect 135594 79778 135622 80036
rect 135686 79898 135714 80036
rect 135778 79937 135806 80036
rect 135764 79928 135820 79937
rect 135674 79892 135726 79898
rect 135764 79863 135820 79872
rect 135674 79834 135726 79840
rect 135870 79812 135898 80036
rect 135306 79766 135358 79772
rect 135456 79750 135622 79778
rect 135718 79792 135774 79801
rect 135352 79416 135404 79422
rect 135352 79358 135404 79364
rect 135168 78056 135220 78062
rect 135168 77998 135220 78004
rect 135076 76492 135128 76498
rect 135076 76434 135128 76440
rect 134984 75472 135036 75478
rect 134984 75414 135036 75420
rect 134708 75268 134760 75274
rect 134708 75210 134760 75216
rect 134628 70366 134748 70394
rect 134720 6662 134748 70366
rect 134708 6656 134760 6662
rect 134708 6598 134760 6604
rect 134524 4140 134576 4146
rect 134524 4082 134576 4088
rect 135364 3602 135392 79358
rect 135456 77926 135484 79750
rect 135718 79727 135774 79736
rect 135824 79784 135898 79812
rect 135628 79688 135680 79694
rect 135628 79630 135680 79636
rect 135536 79552 135588 79558
rect 135536 79494 135588 79500
rect 135548 78033 135576 79494
rect 135534 78024 135590 78033
rect 135534 77959 135590 77968
rect 135444 77920 135496 77926
rect 135444 77862 135496 77868
rect 135640 77518 135668 79630
rect 135628 77512 135680 77518
rect 135628 77454 135680 77460
rect 135628 76832 135680 76838
rect 135628 76774 135680 76780
rect 135444 75336 135496 75342
rect 135444 75278 135496 75284
rect 135456 3738 135484 75278
rect 135536 75200 135588 75206
rect 135536 75142 135588 75148
rect 135548 3874 135576 75142
rect 135536 3868 135588 3874
rect 135536 3810 135588 3816
rect 135444 3732 135496 3738
rect 135444 3674 135496 3680
rect 135640 3670 135668 76774
rect 135732 75914 135760 79727
rect 135824 76838 135852 79784
rect 135962 79744 135990 80036
rect 136054 79971 136082 80036
rect 136040 79962 136096 79971
rect 136040 79897 136096 79906
rect 136146 79898 136174 80036
rect 136134 79892 136186 79898
rect 136134 79834 136186 79840
rect 136238 79744 136266 80036
rect 136330 79898 136358 80036
rect 136422 79898 136450 80036
rect 136318 79892 136370 79898
rect 136318 79834 136370 79840
rect 136410 79892 136462 79898
rect 136410 79834 136462 79840
rect 136514 79830 136542 80036
rect 136606 79966 136634 80036
rect 136594 79960 136646 79966
rect 136594 79902 136646 79908
rect 136502 79824 136554 79830
rect 136698 79812 136726 80036
rect 136790 79830 136818 80036
rect 136882 79830 136910 80036
rect 136974 79898 137002 80036
rect 137066 79898 137094 80036
rect 137158 79971 137186 80036
rect 137144 79962 137200 79971
rect 136962 79892 137014 79898
rect 136962 79834 137014 79840
rect 137054 79892 137106 79898
rect 137144 79897 137200 79906
rect 137250 79898 137278 80036
rect 137342 79971 137370 80036
rect 137328 79962 137384 79971
rect 137434 79966 137462 80036
rect 137526 79966 137554 80036
rect 137618 79966 137646 80036
rect 137710 79966 137738 80036
rect 137054 79834 137106 79840
rect 137238 79892 137290 79898
rect 137328 79897 137384 79906
rect 137422 79960 137474 79966
rect 137422 79902 137474 79908
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137698 79960 137750 79966
rect 137698 79902 137750 79908
rect 137238 79834 137290 79840
rect 136502 79766 136554 79772
rect 136652 79784 136726 79812
rect 136778 79824 136830 79830
rect 135916 79716 135990 79744
rect 136192 79716 136266 79744
rect 135916 77994 135944 79716
rect 136086 79656 136142 79665
rect 136086 79591 136142 79600
rect 135996 79552 136048 79558
rect 135996 79494 136048 79500
rect 135904 77988 135956 77994
rect 135904 77930 135956 77936
rect 135812 76832 135864 76838
rect 135812 76774 135864 76780
rect 135732 75886 135852 75914
rect 135720 75132 135772 75138
rect 135720 75074 135772 75080
rect 135732 11778 135760 75074
rect 135824 11898 135852 75886
rect 135904 75268 135956 75274
rect 135904 75210 135956 75216
rect 135812 11892 135864 11898
rect 135812 11834 135864 11840
rect 135732 11750 135852 11778
rect 135720 11688 135772 11694
rect 135720 11630 135772 11636
rect 135732 3806 135760 11630
rect 135824 4010 135852 11750
rect 135812 4004 135864 4010
rect 135812 3946 135864 3952
rect 135720 3800 135772 3806
rect 135720 3742 135772 3748
rect 135916 3670 135944 75210
rect 136008 45014 136036 79494
rect 135996 45008 136048 45014
rect 135996 44950 136048 44956
rect 136100 6914 136128 79591
rect 136192 75342 136220 79716
rect 136548 79620 136600 79626
rect 136548 79562 136600 79568
rect 136272 79552 136324 79558
rect 136272 79494 136324 79500
rect 136364 79552 136416 79558
rect 136364 79494 136416 79500
rect 136180 75336 136232 75342
rect 136180 75278 136232 75284
rect 136284 75206 136312 79494
rect 136376 75274 136404 79494
rect 136560 78112 136588 79562
rect 136468 78084 136588 78112
rect 136364 75268 136416 75274
rect 136364 75210 136416 75216
rect 136272 75200 136324 75206
rect 136272 75142 136324 75148
rect 136468 75138 136496 78084
rect 136548 77920 136600 77926
rect 136548 77862 136600 77868
rect 136456 75132 136508 75138
rect 136456 75074 136508 75080
rect 136560 75070 136588 77862
rect 136652 77586 136680 79784
rect 136778 79766 136830 79772
rect 136870 79824 136922 79830
rect 137802 79812 137830 80036
rect 136870 79766 136922 79772
rect 137190 79792 137246 79801
rect 137100 79756 137152 79762
rect 137558 79792 137614 79801
rect 137190 79727 137246 79736
rect 137284 79756 137336 79762
rect 137100 79698 137152 79704
rect 136732 79688 136784 79694
rect 136784 79636 136864 79642
rect 136732 79630 136864 79636
rect 136744 79614 136864 79630
rect 136732 79484 136784 79490
rect 136732 79426 136784 79432
rect 136640 77580 136692 77586
rect 136640 77522 136692 77528
rect 136548 75064 136600 75070
rect 136548 75006 136600 75012
rect 136008 6886 136128 6914
rect 135628 3664 135680 3670
rect 135628 3606 135680 3612
rect 135904 3664 135956 3670
rect 135904 3606 135956 3612
rect 135352 3596 135404 3602
rect 135352 3538 135404 3544
rect 136008 3482 136036 6886
rect 136744 3602 136772 79426
rect 136836 75478 136864 79614
rect 136916 79620 136968 79626
rect 136916 79562 136968 79568
rect 136928 77450 136956 79562
rect 137008 79552 137060 79558
rect 137008 79494 137060 79500
rect 136916 77444 136968 77450
rect 136916 77386 136968 77392
rect 136824 75472 136876 75478
rect 136824 75414 136876 75420
rect 136916 75404 136968 75410
rect 136916 75346 136968 75352
rect 136824 75268 136876 75274
rect 136824 75210 136876 75216
rect 136836 3806 136864 75210
rect 136928 4962 136956 75346
rect 137020 75206 137048 79494
rect 137008 75200 137060 75206
rect 137008 75142 137060 75148
rect 137008 75064 137060 75070
rect 137008 75006 137060 75012
rect 136916 4956 136968 4962
rect 136916 4898 136968 4904
rect 137020 4894 137048 75006
rect 137112 5098 137140 79698
rect 137204 75290 137232 79727
rect 137558 79727 137614 79736
rect 137756 79784 137830 79812
rect 137284 79698 137336 79704
rect 137296 75410 137324 79698
rect 137376 79688 137428 79694
rect 137376 79630 137428 79636
rect 137388 76566 137416 79630
rect 137468 79552 137520 79558
rect 137468 79494 137520 79500
rect 137376 76560 137428 76566
rect 137376 76502 137428 76508
rect 137284 75404 137336 75410
rect 137284 75346 137336 75352
rect 137204 75262 137324 75290
rect 137480 75274 137508 79494
rect 137192 75200 137244 75206
rect 137192 75142 137244 75148
rect 137204 60042 137232 75142
rect 137296 66230 137324 75262
rect 137468 75268 137520 75274
rect 137468 75210 137520 75216
rect 137572 73234 137600 79727
rect 137652 75472 137704 75478
rect 137652 75414 137704 75420
rect 137560 73228 137612 73234
rect 137560 73170 137612 73176
rect 137664 70394 137692 75414
rect 137756 75070 137784 79784
rect 137894 79744 137922 80036
rect 137986 79801 138014 80036
rect 138078 79966 138106 80036
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 138170 79898 138198 80036
rect 138262 79898 138290 80036
rect 138158 79892 138210 79898
rect 138158 79834 138210 79840
rect 138250 79892 138302 79898
rect 138250 79834 138302 79840
rect 137848 79716 137922 79744
rect 137972 79792 138028 79801
rect 137972 79727 138028 79736
rect 137848 78169 137876 79716
rect 138020 79688 138072 79694
rect 138354 79676 138382 80036
rect 138446 79971 138474 80036
rect 138432 79962 138488 79971
rect 138538 79966 138566 80036
rect 138630 79966 138658 80036
rect 138432 79897 138488 79906
rect 138526 79960 138578 79966
rect 138526 79902 138578 79908
rect 138618 79960 138670 79966
rect 138618 79902 138670 79908
rect 138722 79744 138750 80036
rect 138814 79778 138842 80036
rect 138906 79898 138934 80036
rect 138998 79937 139026 80036
rect 138984 79928 139040 79937
rect 138894 79892 138946 79898
rect 138984 79863 139040 79872
rect 138894 79834 138946 79840
rect 139090 79830 139118 80036
rect 139078 79824 139130 79830
rect 138814 79750 138934 79778
rect 139182 79801 139210 80036
rect 139274 79966 139302 80036
rect 139366 79966 139394 80036
rect 139458 79966 139486 80036
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139354 79960 139406 79966
rect 139354 79902 139406 79908
rect 139446 79960 139498 79966
rect 139550 79937 139578 80036
rect 139446 79902 139498 79908
rect 139536 79928 139592 79937
rect 139642 79898 139670 80036
rect 139536 79863 139592 79872
rect 139630 79892 139682 79898
rect 139630 79834 139682 79840
rect 139446 79824 139498 79830
rect 139078 79766 139130 79772
rect 139168 79792 139224 79801
rect 138020 79630 138072 79636
rect 138216 79648 138382 79676
rect 138676 79716 138750 79744
rect 137834 78160 137890 78169
rect 137834 78095 137890 78104
rect 138032 78033 138060 79630
rect 138018 78024 138074 78033
rect 138018 77959 138074 77968
rect 138020 77716 138072 77722
rect 138020 77658 138072 77664
rect 137744 75064 137796 75070
rect 137744 75006 137796 75012
rect 137664 70366 137784 70394
rect 137284 66224 137336 66230
rect 137284 66166 137336 66172
rect 137192 60036 137244 60042
rect 137192 59978 137244 59984
rect 137100 5092 137152 5098
rect 137100 5034 137152 5040
rect 137008 4888 137060 4894
rect 137008 4830 137060 4836
rect 137756 3942 137784 70366
rect 138032 5030 138060 77658
rect 138112 75268 138164 75274
rect 138112 75210 138164 75216
rect 138124 5234 138152 75210
rect 138112 5228 138164 5234
rect 138112 5170 138164 5176
rect 138020 5024 138072 5030
rect 138020 4966 138072 4972
rect 138216 4826 138244 79648
rect 138480 79620 138532 79626
rect 138480 79562 138532 79568
rect 138388 79552 138440 79558
rect 138388 79494 138440 79500
rect 138296 79348 138348 79354
rect 138296 79290 138348 79296
rect 138308 6186 138336 79290
rect 138400 20126 138428 79494
rect 138492 44878 138520 79562
rect 138570 78840 138626 78849
rect 138570 78775 138626 78784
rect 138584 66162 138612 78775
rect 138676 75274 138704 79716
rect 138756 79620 138808 79626
rect 138906 79608 138934 79750
rect 139168 79727 139224 79736
rect 139320 79772 139446 79778
rect 139320 79766 139498 79772
rect 139582 79792 139638 79801
rect 139320 79750 139486 79766
rect 138756 79562 138808 79568
rect 138860 79580 138934 79608
rect 139032 79620 139084 79626
rect 138664 75268 138716 75274
rect 138664 75210 138716 75216
rect 138768 75138 138796 79562
rect 138756 75132 138808 75138
rect 138756 75074 138808 75080
rect 138860 70394 138888 79580
rect 139032 79562 139084 79568
rect 139124 79620 139176 79626
rect 139124 79562 139176 79568
rect 138940 79484 138992 79490
rect 138940 79426 138992 79432
rect 138952 71058 138980 79426
rect 139044 77722 139072 79562
rect 139032 77716 139084 77722
rect 139032 77658 139084 77664
rect 139032 77580 139084 77586
rect 139032 77522 139084 77528
rect 138940 71052 138992 71058
rect 138940 70994 138992 71000
rect 138676 70378 138888 70394
rect 138664 70372 138888 70378
rect 138716 70366 138888 70372
rect 138664 70314 138716 70320
rect 138572 66156 138624 66162
rect 138572 66098 138624 66104
rect 139044 64874 139072 77522
rect 139136 75721 139164 79562
rect 139320 77722 139348 79750
rect 139734 79778 139762 80036
rect 139826 79966 139854 80036
rect 139814 79960 139866 79966
rect 139814 79902 139866 79908
rect 139918 79898 139946 80036
rect 140010 79971 140038 80036
rect 139996 79962 140052 79971
rect 140102 79966 140130 80036
rect 139906 79892 139958 79898
rect 139996 79897 140052 79906
rect 140090 79960 140142 79966
rect 140090 79902 140142 79908
rect 139906 79834 139958 79840
rect 139582 79727 139638 79736
rect 139688 79750 139762 79778
rect 139950 79792 140006 79801
rect 139860 79756 139912 79762
rect 139492 79688 139544 79694
rect 139398 79656 139454 79665
rect 139492 79630 139544 79636
rect 139398 79591 139454 79600
rect 139308 77716 139360 77722
rect 139308 77658 139360 77664
rect 139122 75712 139178 75721
rect 139122 75647 139178 75656
rect 138952 64846 139072 64874
rect 138664 60036 138716 60042
rect 138664 59978 138716 59984
rect 138480 44872 138532 44878
rect 138480 44814 138532 44820
rect 138388 20120 138440 20126
rect 138388 20062 138440 20068
rect 138296 6180 138348 6186
rect 138296 6122 138348 6128
rect 138204 4820 138256 4826
rect 138204 4762 138256 4768
rect 138676 4078 138704 59978
rect 138952 4418 138980 64846
rect 139412 27266 139440 79591
rect 139400 27260 139452 27266
rect 139400 27202 139452 27208
rect 139504 27198 139532 79630
rect 139596 28490 139624 79727
rect 139688 78606 139716 79750
rect 140194 79744 140222 80036
rect 140286 79966 140314 80036
rect 140378 79966 140406 80036
rect 140274 79960 140326 79966
rect 140274 79902 140326 79908
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140320 79824 140372 79830
rect 140470 79778 140498 80036
rect 140562 79966 140590 80036
rect 140550 79960 140602 79966
rect 140654 79937 140682 80036
rect 140746 79966 140774 80036
rect 140838 79966 140866 80036
rect 140734 79960 140786 79966
rect 140550 79902 140602 79908
rect 140640 79928 140696 79937
rect 140734 79902 140786 79908
rect 140826 79960 140878 79966
rect 140826 79902 140878 79908
rect 140930 79898 140958 80036
rect 141022 79898 141050 80036
rect 141114 79971 141142 80036
rect 141100 79962 141156 79971
rect 141206 79966 141234 80036
rect 141298 79966 141326 80036
rect 141390 79966 141418 80036
rect 140640 79863 140696 79872
rect 140918 79892 140970 79898
rect 140918 79834 140970 79840
rect 141010 79892 141062 79898
rect 141100 79897 141156 79906
rect 141194 79960 141246 79966
rect 141194 79902 141246 79908
rect 141286 79960 141338 79966
rect 141286 79902 141338 79908
rect 141378 79960 141430 79966
rect 141378 79902 141430 79908
rect 141482 79898 141510 80036
rect 141574 79966 141602 80036
rect 141666 79966 141694 80036
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141654 79960 141706 79966
rect 141654 79902 141706 79908
rect 141010 79834 141062 79840
rect 141470 79892 141522 79898
rect 141470 79834 141522 79840
rect 140320 79766 140372 79772
rect 139950 79727 139952 79736
rect 139860 79698 139912 79704
rect 140004 79727 140006 79736
rect 139952 79698 140004 79704
rect 140148 79716 140222 79744
rect 139768 79552 139820 79558
rect 139768 79494 139820 79500
rect 139676 78600 139728 78606
rect 139676 78542 139728 78548
rect 139676 75268 139728 75274
rect 139676 75210 139728 75216
rect 139688 34134 139716 75210
rect 139780 46238 139808 79494
rect 139872 61538 139900 79698
rect 139950 79656 140006 79665
rect 140006 79614 140084 79642
rect 139950 79591 140006 79600
rect 139952 79484 140004 79490
rect 139952 79426 140004 79432
rect 139964 75585 139992 79426
rect 139950 75576 140006 75585
rect 139950 75511 140006 75520
rect 139952 75200 140004 75206
rect 139952 75142 140004 75148
rect 139964 67454 139992 75142
rect 140056 68678 140084 79614
rect 140148 75274 140176 79716
rect 140228 79620 140280 79626
rect 140228 79562 140280 79568
rect 140136 75268 140188 75274
rect 140136 75210 140188 75216
rect 140240 75206 140268 79562
rect 140332 78062 140360 79766
rect 140424 79750 140498 79778
rect 140688 79756 140740 79762
rect 140320 78056 140372 78062
rect 140320 77998 140372 78004
rect 140424 75857 140452 79750
rect 140688 79698 140740 79704
rect 140780 79756 140832 79762
rect 140780 79698 140832 79704
rect 140596 79688 140648 79694
rect 140596 79630 140648 79636
rect 140504 79416 140556 79422
rect 140504 79358 140556 79364
rect 140410 75848 140466 75857
rect 140410 75783 140466 75792
rect 140228 75200 140280 75206
rect 140228 75142 140280 75148
rect 140412 75132 140464 75138
rect 140412 75074 140464 75080
rect 140044 68672 140096 68678
rect 140044 68614 140096 68620
rect 139952 67448 140004 67454
rect 139952 67390 140004 67396
rect 140044 66224 140096 66230
rect 140044 66166 140096 66172
rect 139860 61532 139912 61538
rect 139860 61474 139912 61480
rect 139768 46232 139820 46238
rect 139768 46174 139820 46180
rect 139676 34128 139728 34134
rect 139676 34070 139728 34076
rect 139584 28484 139636 28490
rect 139584 28426 139636 28432
rect 139492 27192 139544 27198
rect 139492 27134 139544 27140
rect 140056 16574 140084 66166
rect 140056 16546 140176 16574
rect 138940 4412 138992 4418
rect 138940 4354 138992 4360
rect 138664 4072 138716 4078
rect 138664 4014 138716 4020
rect 137744 3936 137796 3942
rect 137744 3878 137796 3884
rect 138848 3868 138900 3874
rect 138848 3810 138900 3816
rect 136824 3800 136876 3806
rect 136824 3742 136876 3748
rect 137652 3732 137704 3738
rect 137652 3674 137704 3680
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 136732 3596 136784 3602
rect 136732 3538 136784 3544
rect 135272 3454 136036 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3538
rect 137664 480 137692 3674
rect 138860 480 138888 3810
rect 140148 3806 140176 16546
rect 140424 6254 140452 75074
rect 140516 27334 140544 79358
rect 140608 75993 140636 79630
rect 140594 75984 140650 75993
rect 140594 75919 140650 75928
rect 140700 74089 140728 79698
rect 140792 78538 140820 79698
rect 141758 79676 141786 80036
rect 141850 79744 141878 80036
rect 141942 79966 141970 80036
rect 142034 79971 142062 80036
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142020 79962 142076 79971
rect 142020 79897 142076 79906
rect 141850 79716 141924 79744
rect 141758 79648 141832 79676
rect 140872 79620 140924 79626
rect 140872 79562 140924 79568
rect 141056 79620 141108 79626
rect 141056 79562 141108 79568
rect 141608 79620 141660 79626
rect 141608 79562 141660 79568
rect 140780 78532 140832 78538
rect 140780 78474 140832 78480
rect 140884 78130 140912 79562
rect 140964 79552 141016 79558
rect 140964 79494 141016 79500
rect 140872 78124 140924 78130
rect 140872 78066 140924 78072
rect 140976 75914 141004 79494
rect 141068 76106 141096 79562
rect 141516 79552 141568 79558
rect 141516 79494 141568 79500
rect 141332 79416 141384 79422
rect 141332 79358 141384 79364
rect 141424 79416 141476 79422
rect 141424 79358 141476 79364
rect 141068 76078 141188 76106
rect 140792 75886 141004 75914
rect 141056 75948 141108 75954
rect 141056 75890 141108 75896
rect 140686 74080 140742 74089
rect 140686 74015 140742 74024
rect 140792 28422 140820 75886
rect 140964 74996 141016 75002
rect 140964 74938 141016 74944
rect 140872 72752 140924 72758
rect 140872 72694 140924 72700
rect 140884 30122 140912 72694
rect 140872 30116 140924 30122
rect 140872 30058 140924 30064
rect 140976 30054 141004 74938
rect 141068 33998 141096 75890
rect 141160 34066 141188 76078
rect 141240 75132 141292 75138
rect 141240 75074 141292 75080
rect 141148 34060 141200 34066
rect 141148 34002 141200 34008
rect 141056 33992 141108 33998
rect 141056 33934 141108 33940
rect 141252 33930 141280 75074
rect 141344 65958 141372 79358
rect 141436 72758 141464 79358
rect 141528 75138 141556 79494
rect 141516 75132 141568 75138
rect 141516 75074 141568 75080
rect 141424 72752 141476 72758
rect 141424 72694 141476 72700
rect 141620 71774 141648 79562
rect 141700 79552 141752 79558
rect 141700 79494 141752 79500
rect 141712 75954 141740 79494
rect 141700 75948 141752 75954
rect 141700 75890 141752 75896
rect 141804 75002 141832 79648
rect 141896 79608 141924 79716
rect 142126 79676 142154 80036
rect 142218 79966 142246 80036
rect 142206 79960 142258 79966
rect 142206 79902 142258 79908
rect 142310 79744 142338 80036
rect 142402 79966 142430 80036
rect 142494 79966 142522 80036
rect 142586 79966 142614 80036
rect 142678 79966 142706 80036
rect 142770 79971 142798 80036
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 142482 79960 142534 79966
rect 142482 79902 142534 79908
rect 142574 79960 142626 79966
rect 142574 79902 142626 79908
rect 142666 79960 142718 79966
rect 142666 79902 142718 79908
rect 142756 79962 142812 79971
rect 142756 79897 142812 79906
rect 142712 79824 142764 79830
rect 142526 79792 142582 79801
rect 142310 79716 142384 79744
rect 142582 79750 142660 79778
rect 142862 79801 142890 80036
rect 142954 79830 142982 80036
rect 143046 79830 143074 80036
rect 143138 79830 143166 80036
rect 143230 79966 143258 80036
rect 143322 79971 143350 80036
rect 143218 79960 143270 79966
rect 143218 79902 143270 79908
rect 143308 79962 143364 79971
rect 143308 79897 143364 79906
rect 142942 79824 142994 79830
rect 142712 79766 142764 79772
rect 142848 79792 142904 79801
rect 142526 79727 142582 79736
rect 142080 79665 142154 79676
rect 142066 79656 142154 79665
rect 141896 79580 142016 79608
rect 142122 79648 142154 79656
rect 142356 79676 142384 79716
rect 142356 79648 142430 79676
rect 142066 79591 142122 79600
rect 142252 79620 142304 79626
rect 141884 79416 141936 79422
rect 141884 79358 141936 79364
rect 141792 74996 141844 75002
rect 141792 74938 141844 74944
rect 141436 71746 141648 71774
rect 141332 65952 141384 65958
rect 141332 65894 141384 65900
rect 141436 65890 141464 71746
rect 141896 70394 141924 79358
rect 141988 74254 142016 79580
rect 142252 79562 142304 79568
rect 142068 79552 142120 79558
rect 142068 79494 142120 79500
rect 142080 79422 142108 79494
rect 142068 79416 142120 79422
rect 142068 79358 142120 79364
rect 142264 78402 142292 79562
rect 142402 79540 142430 79648
rect 142356 79512 142430 79540
rect 142252 78396 142304 78402
rect 142252 78338 142304 78344
rect 142160 75948 142212 75954
rect 142160 75890 142212 75896
rect 141976 74248 142028 74254
rect 141976 74190 142028 74196
rect 141528 70366 141924 70394
rect 141528 70106 141556 70366
rect 141516 70100 141568 70106
rect 141516 70042 141568 70048
rect 141516 66156 141568 66162
rect 141516 66098 141568 66104
rect 141424 65884 141476 65890
rect 141424 65826 141476 65832
rect 141240 33924 141292 33930
rect 141240 33866 141292 33872
rect 140964 30048 141016 30054
rect 140964 29990 141016 29996
rect 140780 28416 140832 28422
rect 140780 28358 140832 28364
rect 140504 27328 140556 27334
rect 140504 27270 140556 27276
rect 140412 6248 140464 6254
rect 140412 6190 140464 6196
rect 141240 4004 141292 4010
rect 141240 3946 141292 3952
rect 140136 3800 140188 3806
rect 140136 3742 140188 3748
rect 140044 3664 140096 3670
rect 140044 3606 140096 3612
rect 140056 480 140084 3606
rect 141252 480 141280 3946
rect 141528 3534 141556 66098
rect 142172 5166 142200 75890
rect 142252 75744 142304 75750
rect 142252 75686 142304 75692
rect 142264 7954 142292 75686
rect 142356 24614 142384 79512
rect 142632 78470 142660 79750
rect 142620 78464 142672 78470
rect 142620 78406 142672 78412
rect 142436 77308 142488 77314
rect 142436 77250 142488 77256
rect 142344 24608 142396 24614
rect 142344 24550 142396 24556
rect 142448 24546 142476 77250
rect 142618 76120 142674 76129
rect 142618 76055 142674 76064
rect 142528 75132 142580 75138
rect 142528 75074 142580 75080
rect 142540 26042 142568 75074
rect 142632 65822 142660 76055
rect 142724 68610 142752 79766
rect 142942 79766 142994 79772
rect 143034 79824 143086 79830
rect 143034 79766 143086 79772
rect 143126 79824 143178 79830
rect 143414 79812 143442 80036
rect 143506 79937 143534 80036
rect 143492 79928 143548 79937
rect 143492 79863 143548 79872
rect 143598 79812 143626 80036
rect 143126 79766 143178 79772
rect 143368 79784 143442 79812
rect 143552 79784 143626 79812
rect 142848 79727 142904 79736
rect 142804 79688 142856 79694
rect 142988 79688 143040 79694
rect 142804 79630 142856 79636
rect 142894 79656 142950 79665
rect 142816 77314 142844 79630
rect 142988 79630 143040 79636
rect 143172 79688 143224 79694
rect 143264 79688 143316 79694
rect 143172 79630 143224 79636
rect 143262 79656 143264 79665
rect 143316 79656 143318 79665
rect 142894 79591 142950 79600
rect 142804 77308 142856 77314
rect 142804 77250 142856 77256
rect 142908 77194 142936 79591
rect 142816 77166 142936 77194
rect 142816 75138 142844 77166
rect 143000 75750 143028 79630
rect 143080 79620 143132 79626
rect 143080 79562 143132 79568
rect 143092 75954 143120 79562
rect 143184 76634 143212 79630
rect 143262 79591 143318 79600
rect 143368 79472 143396 79784
rect 143552 79642 143580 79784
rect 143690 79778 143718 80036
rect 143782 79966 143810 80036
rect 143874 79966 143902 80036
rect 143966 79971 143994 80036
rect 143770 79960 143822 79966
rect 143770 79902 143822 79908
rect 143862 79960 143914 79966
rect 143862 79902 143914 79908
rect 143952 79962 144008 79971
rect 143952 79897 144008 79906
rect 144058 79830 144086 80036
rect 144150 79898 144178 80036
rect 144138 79892 144190 79898
rect 144138 79834 144190 79840
rect 144046 79824 144098 79830
rect 143690 79750 143856 79778
rect 144242 79812 144270 80036
rect 144334 79937 144362 80036
rect 144426 79966 144454 80036
rect 144518 79966 144546 80036
rect 144414 79960 144466 79966
rect 144320 79928 144376 79937
rect 144414 79902 144466 79908
rect 144506 79960 144558 79966
rect 144610 79937 144638 80036
rect 144702 79966 144730 80036
rect 144690 79960 144742 79966
rect 144506 79902 144558 79908
rect 144596 79928 144652 79937
rect 144320 79863 144376 79872
rect 144690 79902 144742 79908
rect 144596 79863 144652 79872
rect 144794 79812 144822 80036
rect 144886 79971 144914 80036
rect 144872 79962 144928 79971
rect 144872 79897 144928 79906
rect 144978 79830 145006 80036
rect 145070 79903 145098 80036
rect 145162 79966 145190 80036
rect 145150 79960 145202 79966
rect 145056 79894 145112 79903
rect 145150 79902 145202 79908
rect 144966 79824 145018 79830
rect 145056 79829 145112 79838
rect 144242 79784 144500 79812
rect 144794 79784 144868 79812
rect 144046 79766 144098 79772
rect 143722 79656 143778 79665
rect 143552 79614 143672 79642
rect 143448 79552 143500 79558
rect 143448 79494 143500 79500
rect 143540 79552 143592 79558
rect 143540 79494 143592 79500
rect 143276 79444 143396 79472
rect 143172 76628 143224 76634
rect 143172 76570 143224 76576
rect 143276 75993 143304 79444
rect 143262 75984 143318 75993
rect 143080 75948 143132 75954
rect 143262 75919 143318 75928
rect 143080 75890 143132 75896
rect 142988 75744 143040 75750
rect 142988 75686 143040 75692
rect 142804 75132 142856 75138
rect 142804 75074 142856 75080
rect 143460 74118 143488 79494
rect 143448 74112 143500 74118
rect 143448 74054 143500 74060
rect 142988 73228 143040 73234
rect 142988 73170 143040 73176
rect 142804 70372 142856 70378
rect 142804 70314 142856 70320
rect 142712 68604 142764 68610
rect 142712 68546 142764 68552
rect 142620 65816 142672 65822
rect 142620 65758 142672 65764
rect 142620 45008 142672 45014
rect 142620 44950 142672 44956
rect 142528 26036 142580 26042
rect 142528 25978 142580 25984
rect 142436 24540 142488 24546
rect 142436 24482 142488 24488
rect 142252 7948 142304 7954
rect 142252 7890 142304 7896
rect 142632 6914 142660 44950
rect 142448 6886 142660 6914
rect 142160 5160 142212 5166
rect 142160 5102 142212 5108
rect 141516 3528 141568 3534
rect 141516 3470 141568 3476
rect 142448 480 142476 6886
rect 142816 3466 142844 70314
rect 143000 3874 143028 73170
rect 143552 7886 143580 79494
rect 143644 77654 143672 79614
rect 143722 79591 143778 79600
rect 143632 77648 143684 77654
rect 143632 77590 143684 77596
rect 143632 76220 143684 76226
rect 143632 76162 143684 76168
rect 143644 12034 143672 76162
rect 143736 14822 143764 79591
rect 143828 76090 143856 79750
rect 143908 79620 143960 79626
rect 143908 79562 143960 79568
rect 144092 79620 144144 79626
rect 144092 79562 144144 79568
rect 144184 79620 144236 79626
rect 144184 79562 144236 79568
rect 144276 79620 144328 79626
rect 144276 79562 144328 79568
rect 143920 76090 143948 79562
rect 144000 79484 144052 79490
rect 144000 79426 144052 79432
rect 144012 78878 144040 79426
rect 144000 78872 144052 78878
rect 144000 78814 144052 78820
rect 144104 76226 144132 79562
rect 144092 76220 144144 76226
rect 144092 76162 144144 76168
rect 143816 76084 143868 76090
rect 143816 76026 143868 76032
rect 143908 76084 143960 76090
rect 143908 76026 143960 76032
rect 144092 76084 144144 76090
rect 144092 76026 144144 76032
rect 143814 75984 143870 75993
rect 143814 75919 143870 75928
rect 143908 75948 143960 75954
rect 143828 29918 143856 75919
rect 143908 75890 143960 75896
rect 143920 29986 143948 75890
rect 144000 75268 144052 75274
rect 144000 75210 144052 75216
rect 144012 31482 144040 75210
rect 144104 33862 144132 76026
rect 144196 64462 144224 79562
rect 144288 64530 144316 79562
rect 144472 78946 144500 79784
rect 144552 79756 144604 79762
rect 144552 79698 144604 79704
rect 144644 79756 144696 79762
rect 144840 79744 144868 79784
rect 145254 79812 145282 80036
rect 144966 79766 145018 79772
rect 145208 79784 145282 79812
rect 144644 79698 144696 79704
rect 144748 79716 144868 79744
rect 144460 78940 144512 78946
rect 144460 78882 144512 78888
rect 144564 78826 144592 79698
rect 144472 78798 144592 78826
rect 144472 75274 144500 78798
rect 144656 78713 144684 79698
rect 144642 78704 144698 78713
rect 144642 78639 144698 78648
rect 144748 76945 144776 79716
rect 144920 79688 144972 79694
rect 144920 79630 144972 79636
rect 145012 79688 145064 79694
rect 145012 79630 145064 79636
rect 145102 79656 145158 79665
rect 144828 79620 144880 79626
rect 144828 79562 144880 79568
rect 144734 76936 144790 76945
rect 144734 76871 144790 76880
rect 144552 76560 144604 76566
rect 144552 76502 144604 76508
rect 144460 75268 144512 75274
rect 144460 75210 144512 75216
rect 144564 70394 144592 76502
rect 144840 74186 144868 79562
rect 144932 77382 144960 79630
rect 144920 77376 144972 77382
rect 144920 77318 144972 77324
rect 144920 75336 144972 75342
rect 144920 75278 144972 75284
rect 144828 74180 144880 74186
rect 144828 74122 144880 74128
rect 144472 70366 144592 70394
rect 144276 64524 144328 64530
rect 144276 64466 144328 64472
rect 144184 64456 144236 64462
rect 144184 64398 144236 64404
rect 144092 33856 144144 33862
rect 144092 33798 144144 33804
rect 144000 31476 144052 31482
rect 144000 31418 144052 31424
rect 143908 29980 143960 29986
rect 143908 29922 143960 29928
rect 143816 29912 143868 29918
rect 143816 29854 143868 29860
rect 143724 14816 143776 14822
rect 143724 14758 143776 14764
rect 143632 12028 143684 12034
rect 143632 11970 143684 11976
rect 143540 7880 143592 7886
rect 143540 7822 143592 7828
rect 143540 4412 143592 4418
rect 143540 4354 143592 4360
rect 142988 3868 143040 3874
rect 142988 3810 143040 3816
rect 142804 3460 142856 3466
rect 142804 3402 142856 3408
rect 143552 480 143580 4354
rect 144472 3330 144500 70366
rect 144932 9314 144960 75278
rect 145024 20398 145052 79630
rect 145102 79591 145158 79600
rect 145116 75206 145144 79591
rect 145208 79082 145236 79784
rect 145346 79676 145374 80036
rect 145438 79966 145466 80036
rect 145426 79960 145478 79966
rect 145530 79937 145558 80036
rect 145426 79902 145478 79908
rect 145516 79928 145572 79937
rect 145622 79898 145650 80036
rect 145516 79863 145572 79872
rect 145610 79892 145662 79898
rect 145610 79834 145662 79840
rect 145714 79812 145742 80036
rect 145806 79966 145834 80036
rect 145898 79966 145926 80036
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145886 79960 145938 79966
rect 145990 79937 146018 80036
rect 145886 79902 145938 79908
rect 145976 79928 146032 79937
rect 145976 79863 146032 79872
rect 145840 79824 145892 79830
rect 145714 79784 145788 79812
rect 145300 79648 145374 79676
rect 145656 79688 145708 79694
rect 145470 79656 145526 79665
rect 145196 79076 145248 79082
rect 145196 79018 145248 79024
rect 145196 78872 145248 78878
rect 145196 78814 145248 78820
rect 145104 75200 145156 75206
rect 145104 75142 145156 75148
rect 145104 75064 145156 75070
rect 145104 75006 145156 75012
rect 145012 20392 145064 20398
rect 145012 20334 145064 20340
rect 145116 20330 145144 75006
rect 145208 29782 145236 78814
rect 145300 29850 145328 79648
rect 145656 79630 145708 79636
rect 145470 79591 145526 79600
rect 145380 79552 145432 79558
rect 145380 79494 145432 79500
rect 145392 77294 145420 79494
rect 145484 78656 145512 79591
rect 145668 78878 145696 79630
rect 145656 78872 145708 78878
rect 145656 78814 145708 78820
rect 145656 78668 145708 78674
rect 145484 78628 145604 78656
rect 145392 77266 145512 77294
rect 145484 76702 145512 77266
rect 145472 76696 145524 76702
rect 145472 76638 145524 76644
rect 145380 75268 145432 75274
rect 145380 75210 145432 75216
rect 145392 35630 145420 75210
rect 145472 75200 145524 75206
rect 145472 75142 145524 75148
rect 145484 65754 145512 75142
rect 145472 65748 145524 65754
rect 145472 65690 145524 65696
rect 145576 65686 145604 78628
rect 145656 78610 145708 78616
rect 145668 76838 145696 78610
rect 145656 76832 145708 76838
rect 145656 76774 145708 76780
rect 145656 76696 145708 76702
rect 145656 76638 145708 76644
rect 145668 74050 145696 76638
rect 145760 75274 145788 79784
rect 145840 79766 145892 79772
rect 145852 75342 145880 79766
rect 146082 79744 146110 80036
rect 146174 79937 146202 80036
rect 146160 79928 146216 79937
rect 146160 79863 146216 79872
rect 146082 79716 146156 79744
rect 146024 79552 146076 79558
rect 146024 79494 146076 79500
rect 145930 78840 145986 78849
rect 145930 78775 145986 78784
rect 145840 75336 145892 75342
rect 145840 75278 145892 75284
rect 145748 75268 145800 75274
rect 145748 75210 145800 75216
rect 145944 75070 145972 78775
rect 146036 78674 146064 79494
rect 146024 78668 146076 78674
rect 146024 78610 146076 78616
rect 146128 78577 146156 79716
rect 146266 79676 146294 80036
rect 146358 79937 146386 80036
rect 146344 79928 146400 79937
rect 146344 79863 146400 79872
rect 146450 79744 146478 80036
rect 146220 79648 146294 79676
rect 146404 79716 146478 79744
rect 146220 78713 146248 79648
rect 146300 79552 146352 79558
rect 146300 79494 146352 79500
rect 146206 78704 146262 78713
rect 146206 78639 146262 78648
rect 146114 78568 146170 78577
rect 146114 78503 146170 78512
rect 146208 75336 146260 75342
rect 146208 75278 146260 75284
rect 145932 75064 145984 75070
rect 145932 75006 145984 75012
rect 146220 74746 146248 75278
rect 146312 74934 146340 79494
rect 146404 78928 146432 79716
rect 146542 79608 146570 80036
rect 146634 79830 146662 80036
rect 146622 79824 146674 79830
rect 146622 79766 146674 79772
rect 146726 79676 146754 80036
rect 146680 79648 146754 79676
rect 146542 79580 146616 79608
rect 146404 78900 146524 78928
rect 146392 78668 146444 78674
rect 146392 78610 146444 78616
rect 146300 74928 146352 74934
rect 146300 74870 146352 74876
rect 146220 74718 146340 74746
rect 145656 74044 145708 74050
rect 145656 73986 145708 73992
rect 145564 65680 145616 65686
rect 145564 65622 145616 65628
rect 145380 35624 145432 35630
rect 145380 35566 145432 35572
rect 145288 29844 145340 29850
rect 145288 29786 145340 29792
rect 145196 29776 145248 29782
rect 145196 29718 145248 29724
rect 145104 20324 145156 20330
rect 145104 20266 145156 20272
rect 144920 9308 144972 9314
rect 144920 9250 144972 9256
rect 146312 9246 146340 74718
rect 146404 20262 146432 78610
rect 146496 75274 146524 78900
rect 146484 75268 146536 75274
rect 146484 75210 146536 75216
rect 146588 75206 146616 79580
rect 146576 75200 146628 75206
rect 146576 75142 146628 75148
rect 146484 75132 146536 75138
rect 146484 75074 146536 75080
rect 146496 25974 146524 75074
rect 146576 75064 146628 75070
rect 146576 75006 146628 75012
rect 146588 27130 146616 75006
rect 146680 28354 146708 79648
rect 146818 79608 146846 80036
rect 146910 79778 146938 80036
rect 147002 79898 147030 80036
rect 147094 79966 147122 80036
rect 147082 79960 147134 79966
rect 147082 79902 147134 79908
rect 146990 79892 147042 79898
rect 146990 79834 147042 79840
rect 147186 79778 147214 80036
rect 147278 79898 147306 80036
rect 147370 79971 147398 80036
rect 147356 79962 147412 79971
rect 147462 79966 147490 80036
rect 147266 79892 147318 79898
rect 147356 79897 147412 79906
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147266 79834 147318 79840
rect 147404 79824 147456 79830
rect 146910 79750 147076 79778
rect 147186 79750 147306 79778
rect 147404 79766 147456 79772
rect 146772 79580 146846 79608
rect 146772 78674 146800 79580
rect 146944 79416 146996 79422
rect 146944 79358 146996 79364
rect 146956 79218 146984 79358
rect 146944 79212 146996 79218
rect 146944 79154 146996 79160
rect 146944 78940 146996 78946
rect 146944 78882 146996 78888
rect 146852 78736 146904 78742
rect 146852 78678 146904 78684
rect 146760 78668 146812 78674
rect 146760 78610 146812 78616
rect 146864 75342 146892 78678
rect 146956 76906 146984 78882
rect 146944 76900 146996 76906
rect 146944 76842 146996 76848
rect 146852 75336 146904 75342
rect 146852 75278 146904 75284
rect 146760 75268 146812 75274
rect 146760 75210 146812 75216
rect 146944 75268 146996 75274
rect 146944 75210 146996 75216
rect 146772 31414 146800 75210
rect 146852 75200 146904 75206
rect 146852 75142 146904 75148
rect 146864 33794 146892 75142
rect 146956 35562 146984 75210
rect 147048 63170 147076 79750
rect 147278 79744 147306 79750
rect 147278 79716 147352 79744
rect 147128 79688 147180 79694
rect 147128 79630 147180 79636
rect 147140 75274 147168 79630
rect 147220 79620 147272 79626
rect 147220 79562 147272 79568
rect 147128 75268 147180 75274
rect 147128 75210 147180 75216
rect 147232 75070 147260 79562
rect 147324 78742 147352 79716
rect 147312 78736 147364 78742
rect 147416 78713 147444 79766
rect 147554 79676 147582 80036
rect 147646 79835 147674 80036
rect 147632 79826 147688 79835
rect 147738 79830 147766 80036
rect 147830 79830 147858 80036
rect 147922 79898 147950 80036
rect 148014 79937 148042 80036
rect 148106 79966 148134 80036
rect 148198 79966 148226 80036
rect 148290 79966 148318 80036
rect 148094 79960 148146 79966
rect 148000 79928 148056 79937
rect 147910 79892 147962 79898
rect 148094 79902 148146 79908
rect 148186 79960 148238 79966
rect 148186 79902 148238 79908
rect 148278 79960 148330 79966
rect 148278 79902 148330 79908
rect 148382 79898 148410 80036
rect 148000 79863 148056 79872
rect 148370 79892 148422 79898
rect 147910 79834 147962 79840
rect 148370 79834 148422 79840
rect 147632 79761 147688 79770
rect 147726 79824 147778 79830
rect 147726 79766 147778 79772
rect 147818 79824 147870 79830
rect 148278 79824 148330 79830
rect 147818 79766 147870 79772
rect 148198 79772 148278 79778
rect 148198 79766 148330 79772
rect 147956 79756 148008 79762
rect 147956 79698 148008 79704
rect 148048 79756 148100 79762
rect 148048 79698 148100 79704
rect 148198 79750 148318 79766
rect 147864 79688 147916 79694
rect 147554 79648 147720 79676
rect 147496 79552 147548 79558
rect 147496 79494 147548 79500
rect 147312 78678 147364 78684
rect 147402 78704 147458 78713
rect 147402 78639 147458 78648
rect 147508 75138 147536 79494
rect 147588 79076 147640 79082
rect 147588 79018 147640 79024
rect 147600 78674 147628 79018
rect 147588 78668 147640 78674
rect 147588 78610 147640 78616
rect 147692 76809 147720 79648
rect 147864 79630 147916 79636
rect 147772 79620 147824 79626
rect 147772 79562 147824 79568
rect 147784 77518 147812 79562
rect 147772 77512 147824 77518
rect 147772 77454 147824 77460
rect 147678 76800 147734 76809
rect 147678 76735 147734 76744
rect 147680 75336 147732 75342
rect 147680 75278 147732 75284
rect 147496 75132 147548 75138
rect 147496 75074 147548 75080
rect 147220 75064 147272 75070
rect 147220 75006 147272 75012
rect 147220 74928 147272 74934
rect 147220 74870 147272 74876
rect 147232 67386 147260 74870
rect 147220 67380 147272 67386
rect 147220 67322 147272 67328
rect 147036 63164 147088 63170
rect 147036 63106 147088 63112
rect 147036 44872 147088 44878
rect 147036 44814 147088 44820
rect 146944 35556 146996 35562
rect 146944 35498 146996 35504
rect 146852 33788 146904 33794
rect 146852 33730 146904 33736
rect 146760 31408 146812 31414
rect 146760 31350 146812 31356
rect 146668 28348 146720 28354
rect 146668 28290 146720 28296
rect 146576 27124 146628 27130
rect 146576 27066 146628 27072
rect 146484 25968 146536 25974
rect 146484 25910 146536 25916
rect 146392 20256 146444 20262
rect 146392 20198 146444 20204
rect 147048 16574 147076 44814
rect 147048 16546 147260 16574
rect 146300 9240 146352 9246
rect 146300 9182 146352 9188
rect 145932 4072 145984 4078
rect 145932 4014 145984 4020
rect 144736 3936 144788 3942
rect 144736 3878 144788 3884
rect 144460 3324 144512 3330
rect 144460 3266 144512 3272
rect 144748 480 144776 3878
rect 145944 480 145972 4014
rect 147232 3602 147260 16546
rect 147692 10606 147720 75278
rect 147772 75200 147824 75206
rect 147772 75142 147824 75148
rect 147784 24478 147812 75142
rect 147876 28286 147904 79630
rect 147968 78742 147996 79698
rect 147956 78736 148008 78742
rect 147956 78678 148008 78684
rect 148060 77294 148088 79698
rect 148198 79676 148226 79750
rect 148474 79744 148502 80036
rect 148428 79716 148502 79744
rect 148324 79688 148376 79694
rect 148198 79648 148272 79676
rect 148140 78736 148192 78742
rect 148140 78678 148192 78684
rect 147968 77266 148088 77294
rect 147968 31346 147996 77266
rect 148048 75268 148100 75274
rect 148048 75210 148100 75216
rect 148060 35426 148088 75210
rect 148152 35494 148180 78678
rect 148244 64394 148272 79648
rect 148324 79630 148376 79636
rect 148336 78878 148364 79630
rect 148324 78872 148376 78878
rect 148324 78814 148376 78820
rect 148324 78736 148376 78742
rect 148324 78678 148376 78684
rect 148336 76770 148364 78678
rect 148324 76764 148376 76770
rect 148324 76706 148376 76712
rect 148428 75274 148456 79716
rect 148566 79608 148594 80036
rect 148658 79676 148686 80036
rect 148750 79937 148778 80036
rect 148736 79928 148792 79937
rect 148842 79898 148870 80036
rect 148736 79863 148792 79872
rect 148830 79892 148882 79898
rect 148830 79834 148882 79840
rect 148934 79801 148962 80036
rect 149026 79966 149054 80036
rect 149118 79966 149146 80036
rect 149014 79960 149066 79966
rect 149014 79902 149066 79908
rect 149106 79960 149158 79966
rect 149106 79902 149158 79908
rect 148920 79792 148976 79801
rect 148784 79756 148836 79762
rect 149210 79778 149238 80036
rect 148920 79727 148976 79736
rect 149164 79750 149238 79778
rect 149302 79778 149330 80036
rect 149394 79898 149422 80036
rect 149486 79966 149514 80036
rect 149474 79960 149526 79966
rect 149474 79902 149526 79908
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 149578 79778 149606 80036
rect 149302 79750 149376 79778
rect 148784 79698 148836 79704
rect 148658 79648 148732 79676
rect 148566 79580 148640 79608
rect 148508 78872 148560 78878
rect 148508 78814 148560 78820
rect 148416 75268 148468 75274
rect 148416 75210 148468 75216
rect 148520 75206 148548 78814
rect 148612 75342 148640 79580
rect 148704 78742 148732 79648
rect 148692 78736 148744 78742
rect 148796 78713 148824 79698
rect 149060 79688 149112 79694
rect 148966 79656 149022 79665
rect 148876 79620 148928 79626
rect 149060 79630 149112 79636
rect 148966 79591 149022 79600
rect 148876 79562 148928 79568
rect 148692 78678 148744 78684
rect 148782 78704 148838 78713
rect 148782 78639 148838 78648
rect 148888 78441 148916 79562
rect 148980 79082 149008 79591
rect 148968 79076 149020 79082
rect 148968 79018 149020 79024
rect 149072 78849 149100 79630
rect 149058 78840 149114 78849
rect 149058 78775 149114 78784
rect 149058 78704 149114 78713
rect 149058 78639 149114 78648
rect 148874 78432 148930 78441
rect 148874 78367 148930 78376
rect 148692 78056 148744 78062
rect 148692 77998 148744 78004
rect 148600 75336 148652 75342
rect 148600 75278 148652 75284
rect 148508 75200 148560 75206
rect 148508 75142 148560 75148
rect 148232 64388 148284 64394
rect 148232 64330 148284 64336
rect 148140 35488 148192 35494
rect 148140 35430 148192 35436
rect 148048 35420 148100 35426
rect 148048 35362 148100 35368
rect 147956 31340 148008 31346
rect 147956 31282 148008 31288
rect 148704 28558 148732 77998
rect 148874 77480 148930 77489
rect 148874 77415 148930 77424
rect 148888 77314 148916 77415
rect 148876 77308 148928 77314
rect 148876 77250 148928 77256
rect 148968 77240 149020 77246
rect 148968 77182 149020 77188
rect 148980 72690 149008 77182
rect 148968 72684 149020 72690
rect 148968 72626 149020 72632
rect 149072 72622 149100 78639
rect 149060 72616 149112 72622
rect 149060 72558 149112 72564
rect 148692 28552 148744 28558
rect 148692 28494 148744 28500
rect 147864 28280 147916 28286
rect 147864 28222 147916 28228
rect 147772 24472 147824 24478
rect 147772 24414 147824 24420
rect 149164 23390 149192 79750
rect 149244 79688 149296 79694
rect 149244 79630 149296 79636
rect 149256 25906 149284 79630
rect 149348 75410 149376 79750
rect 149532 79750 149606 79778
rect 149532 79676 149560 79750
rect 149670 79676 149698 80036
rect 149762 79966 149790 80036
rect 149750 79960 149802 79966
rect 149854 79937 149882 80036
rect 149750 79902 149802 79908
rect 149840 79928 149896 79937
rect 149840 79863 149896 79872
rect 149946 79812 149974 80036
rect 150038 79966 150066 80036
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 150130 79898 150158 80036
rect 150222 79903 150250 80036
rect 150118 79892 150170 79898
rect 150118 79834 150170 79840
rect 150208 79894 150264 79903
rect 150208 79829 150264 79838
rect 149946 79784 150066 79812
rect 149440 79648 149560 79676
rect 149624 79648 149698 79676
rect 149796 79688 149848 79694
rect 149336 75404 149388 75410
rect 149336 75346 149388 75352
rect 149336 75268 149388 75274
rect 149336 75210 149388 75216
rect 149348 27062 149376 75210
rect 149440 35290 149468 79648
rect 149520 79552 149572 79558
rect 149520 79494 149572 79500
rect 149532 77246 149560 79494
rect 149520 77240 149572 77246
rect 149520 77182 149572 77188
rect 149520 75404 149572 75410
rect 149520 75346 149572 75352
rect 149532 35358 149560 75346
rect 149624 63102 149652 79648
rect 150038 79676 150066 79784
rect 150164 79756 150216 79762
rect 150314 79744 150342 80036
rect 150406 79903 150434 80036
rect 150498 79966 150526 80036
rect 150486 79960 150538 79966
rect 150392 79894 150448 79903
rect 150486 79902 150538 79908
rect 150392 79829 150448 79838
rect 150164 79698 150216 79704
rect 150268 79716 150342 79744
rect 150590 79744 150618 80036
rect 150682 79812 150710 80036
rect 150774 79966 150802 80036
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150682 79784 150756 79812
rect 150866 79801 150894 80036
rect 150958 79830 150986 80036
rect 151050 79937 151078 80036
rect 151036 79928 151092 79937
rect 151036 79863 151092 79872
rect 150946 79824 150998 79830
rect 150590 79716 150664 79744
rect 150038 79648 150112 79676
rect 149796 79630 149848 79636
rect 149704 79416 149756 79422
rect 149704 79358 149756 79364
rect 149716 79218 149744 79358
rect 149704 79212 149756 79218
rect 149704 79154 149756 79160
rect 149702 78840 149758 78849
rect 149702 78775 149758 78784
rect 149716 77450 149744 78775
rect 149704 77444 149756 77450
rect 149704 77386 149756 77392
rect 149808 70394 149836 79630
rect 149888 79620 149940 79626
rect 149888 79562 149940 79568
rect 149900 75274 149928 79562
rect 150084 78418 150112 79648
rect 150176 78577 150204 79698
rect 150268 78713 150296 79716
rect 150348 79620 150400 79626
rect 150400 79580 150572 79608
rect 150348 79562 150400 79568
rect 150348 79280 150400 79286
rect 150348 79222 150400 79228
rect 150360 79150 150388 79222
rect 150348 79144 150400 79150
rect 150348 79086 150400 79092
rect 150254 78704 150310 78713
rect 150254 78639 150310 78648
rect 150438 78704 150494 78713
rect 150438 78639 150494 78648
rect 150162 78568 150218 78577
rect 150162 78503 150218 78512
rect 150084 78390 150388 78418
rect 150256 78056 150308 78062
rect 150256 77998 150308 78004
rect 150268 76498 150296 77998
rect 150256 76492 150308 76498
rect 150256 76434 150308 76440
rect 149888 75268 149940 75274
rect 149888 75210 149940 75216
rect 149716 70366 149836 70394
rect 149716 67318 149744 70366
rect 149704 67312 149756 67318
rect 149704 67254 149756 67260
rect 149612 63096 149664 63102
rect 149612 63038 149664 63044
rect 149520 35352 149572 35358
rect 149520 35294 149572 35300
rect 149428 35284 149480 35290
rect 149428 35226 149480 35232
rect 149336 27056 149388 27062
rect 149336 26998 149388 27004
rect 149244 25900 149296 25906
rect 149244 25842 149296 25848
rect 149152 23384 149204 23390
rect 149152 23326 149204 23332
rect 150360 11966 150388 78390
rect 150452 70394 150480 78639
rect 150544 76702 150572 79580
rect 150532 76696 150584 76702
rect 150532 76638 150584 76644
rect 150452 70366 150572 70394
rect 150348 11960 150400 11966
rect 150348 11902 150400 11908
rect 147680 10600 147732 10606
rect 147680 10542 147732 10548
rect 148324 5092 148376 5098
rect 148324 5034 148376 5040
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 147220 3596 147272 3602
rect 147220 3538 147272 3544
rect 147140 480 147168 3538
rect 148336 480 148364 5034
rect 150544 4078 150572 70366
rect 150636 5114 150664 79716
rect 150728 75274 150756 79784
rect 150852 79792 150908 79801
rect 150946 79766 150998 79772
rect 151142 79744 151170 80036
rect 151234 79966 151262 80036
rect 151326 79971 151354 80036
rect 151222 79960 151274 79966
rect 151222 79902 151274 79908
rect 151312 79962 151368 79971
rect 151312 79897 151368 79906
rect 151418 79744 151446 80036
rect 151510 79966 151538 80036
rect 151602 79966 151630 80036
rect 151694 79966 151722 80036
rect 151498 79960 151550 79966
rect 151498 79902 151550 79908
rect 151590 79960 151642 79966
rect 151590 79902 151642 79908
rect 151682 79960 151734 79966
rect 151786 79937 151814 80036
rect 151682 79902 151734 79908
rect 151772 79928 151828 79937
rect 151878 79898 151906 80036
rect 151970 79966 151998 80036
rect 152062 79966 152090 80036
rect 152154 79966 152182 80036
rect 152246 79971 152274 80036
rect 151958 79960 152010 79966
rect 151958 79902 152010 79908
rect 152050 79960 152102 79966
rect 152050 79902 152102 79908
rect 152142 79960 152194 79966
rect 152142 79902 152194 79908
rect 152232 79962 152288 79971
rect 151772 79863 151828 79872
rect 151866 79892 151918 79898
rect 152232 79897 152288 79906
rect 151866 79834 151918 79840
rect 150852 79727 150908 79736
rect 151096 79716 151170 79744
rect 151372 79716 151446 79744
rect 151726 79792 151782 79801
rect 152186 79792 152242 79801
rect 151726 79727 151782 79736
rect 151820 79756 151872 79762
rect 150808 79688 150860 79694
rect 150808 79630 150860 79636
rect 150900 79688 150952 79694
rect 150900 79630 150952 79636
rect 150992 79688 151044 79694
rect 150992 79630 151044 79636
rect 150716 75268 150768 75274
rect 150716 75210 150768 75216
rect 150716 75132 150768 75138
rect 150716 75074 150768 75080
rect 150728 5386 150756 75074
rect 150820 6594 150848 79630
rect 150912 6730 150940 79630
rect 151004 77897 151032 79630
rect 150990 77888 151046 77897
rect 150990 77823 151046 77832
rect 151096 77294 151124 79716
rect 151372 79676 151400 79716
rect 151326 79648 151400 79676
rect 151176 79620 151228 79626
rect 151176 79562 151228 79568
rect 151188 78713 151216 79562
rect 151326 79540 151354 79648
rect 151740 79642 151768 79727
rect 152338 79778 152366 80036
rect 152430 79971 152458 80036
rect 152416 79962 152472 79971
rect 152522 79966 152550 80036
rect 152416 79897 152472 79906
rect 152510 79960 152562 79966
rect 152614 79937 152642 80036
rect 152510 79902 152562 79908
rect 152600 79928 152656 79937
rect 152706 79898 152734 80036
rect 152600 79863 152656 79872
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 152186 79727 152242 79736
rect 152292 79750 152366 79778
rect 152556 79824 152608 79830
rect 152556 79766 152608 79772
rect 152646 79792 152702 79801
rect 151820 79698 151872 79704
rect 151648 79614 151768 79642
rect 151280 79512 151354 79540
rect 151544 79552 151596 79558
rect 151174 78704 151230 78713
rect 151174 78639 151230 78648
rect 151280 77314 151308 79512
rect 151544 79494 151596 79500
rect 151452 79484 151504 79490
rect 151452 79426 151504 79432
rect 151464 79150 151492 79426
rect 151452 79144 151504 79150
rect 151452 79086 151504 79092
rect 151358 78840 151414 78849
rect 151358 78775 151414 78784
rect 151004 77266 151124 77294
rect 151268 77308 151320 77314
rect 150900 6724 150952 6730
rect 150900 6666 150952 6672
rect 151004 6662 151032 77266
rect 151268 77250 151320 77256
rect 151084 75268 151136 75274
rect 151084 75210 151136 75216
rect 151096 6798 151124 75210
rect 151372 75138 151400 78775
rect 151556 77858 151584 79494
rect 151544 77852 151596 77858
rect 151544 77794 151596 77800
rect 151648 77294 151676 79614
rect 151728 79552 151780 79558
rect 151728 79494 151780 79500
rect 151740 78577 151768 79494
rect 151726 78568 151782 78577
rect 151726 78503 151782 78512
rect 151464 77266 151676 77294
rect 151360 75132 151412 75138
rect 151360 75074 151412 75080
rect 151464 70394 151492 77266
rect 151832 76294 151860 79698
rect 152002 79656 152058 79665
rect 151912 79620 151964 79626
rect 152002 79591 152058 79600
rect 151912 79562 151964 79568
rect 151820 76288 151872 76294
rect 151820 76230 151872 76236
rect 151820 75744 151872 75750
rect 151820 75686 151872 75692
rect 151464 70366 151584 70394
rect 151084 6792 151136 6798
rect 151084 6734 151136 6740
rect 150992 6656 151044 6662
rect 150992 6598 151044 6604
rect 150808 6588 150860 6594
rect 150808 6530 150860 6536
rect 150728 5358 150940 5386
rect 150636 5086 150848 5114
rect 150624 4956 150676 4962
rect 150624 4898 150676 4904
rect 150532 4072 150584 4078
rect 150532 4014 150584 4020
rect 149520 3800 149572 3806
rect 149520 3742 149572 3748
rect 149532 480 149560 3742
rect 150636 480 150664 4898
rect 150820 3398 150848 5086
rect 150912 4010 150940 5358
rect 151556 4146 151584 70366
rect 151832 9178 151860 75686
rect 151924 75342 151952 79562
rect 151912 75336 151964 75342
rect 151912 75278 151964 75284
rect 151912 75200 151964 75206
rect 151912 75142 151964 75148
rect 151924 13394 151952 75142
rect 152016 13462 152044 79591
rect 152096 76560 152148 76566
rect 152096 76502 152148 76508
rect 152108 21690 152136 76502
rect 152200 75750 152228 79727
rect 152292 76566 152320 79750
rect 152464 79620 152516 79626
rect 152464 79562 152516 79568
rect 152372 76968 152424 76974
rect 152372 76910 152424 76916
rect 152384 76634 152412 76910
rect 152372 76628 152424 76634
rect 152372 76570 152424 76576
rect 152280 76560 152332 76566
rect 152280 76502 152332 76508
rect 152280 76288 152332 76294
rect 152280 76230 152332 76236
rect 152188 75744 152240 75750
rect 152188 75686 152240 75692
rect 152188 75268 152240 75274
rect 152188 75210 152240 75216
rect 152200 25838 152228 75210
rect 152292 26994 152320 76230
rect 152372 75336 152424 75342
rect 152372 75278 152424 75284
rect 152384 64326 152412 75278
rect 152476 67182 152504 79562
rect 152568 75274 152596 79766
rect 152646 79727 152702 79736
rect 152798 79744 152826 80036
rect 152890 79937 152918 80036
rect 152982 79966 153010 80036
rect 152970 79960 153022 79966
rect 152876 79928 152932 79937
rect 152970 79902 153022 79908
rect 152876 79863 152932 79872
rect 153074 79812 153102 80036
rect 153166 79971 153194 80036
rect 153152 79962 153208 79971
rect 153258 79966 153286 80036
rect 153152 79897 153208 79906
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153028 79801 153102 79812
rect 153014 79792 153102 79801
rect 152660 78334 152688 79727
rect 152798 79716 152872 79744
rect 153070 79784 153102 79792
rect 153350 79744 153378 80036
rect 153014 79727 153070 79736
rect 152740 79552 152792 79558
rect 152740 79494 152792 79500
rect 152648 78328 152700 78334
rect 152648 78270 152700 78276
rect 152648 77444 152700 77450
rect 152648 77386 152700 77392
rect 152556 75268 152608 75274
rect 152556 75210 152608 75216
rect 152660 73982 152688 77386
rect 152648 73976 152700 73982
rect 152648 73918 152700 73924
rect 152752 72554 152780 79494
rect 152844 76673 152872 79716
rect 153212 79716 153378 79744
rect 153016 79688 153068 79694
rect 153016 79630 153068 79636
rect 153106 79656 153162 79665
rect 152924 79620 152976 79626
rect 152924 79562 152976 79568
rect 152830 76664 152886 76673
rect 152830 76599 152886 76608
rect 152936 75206 152964 79562
rect 153028 77353 153056 79630
rect 153106 79591 153162 79600
rect 153014 77344 153070 77353
rect 153014 77279 153070 77288
rect 153016 77240 153068 77246
rect 153016 77182 153068 77188
rect 153028 76770 153056 77182
rect 153016 76764 153068 76770
rect 153016 76706 153068 76712
rect 152924 75200 152976 75206
rect 152924 75142 152976 75148
rect 153120 73914 153148 79591
rect 153212 76106 153240 79716
rect 153442 79676 153470 80036
rect 153534 79830 153562 80036
rect 153626 79966 153654 80036
rect 153614 79960 153666 79966
rect 153614 79902 153666 79908
rect 153718 79898 153746 80036
rect 153810 79966 153838 80036
rect 153902 79971 153930 80036
rect 153798 79960 153850 79966
rect 153798 79902 153850 79908
rect 153888 79962 153944 79971
rect 153706 79892 153758 79898
rect 153888 79897 153944 79906
rect 153706 79834 153758 79840
rect 153522 79824 153574 79830
rect 153522 79766 153574 79772
rect 153994 79778 154022 80036
rect 154086 79966 154114 80036
rect 154074 79960 154126 79966
rect 154074 79902 154126 79908
rect 154178 79830 154206 80036
rect 154166 79824 154218 79830
rect 153660 79756 153712 79762
rect 153994 79750 154068 79778
rect 154166 79766 154218 79772
rect 153660 79698 153712 79704
rect 153568 79688 153620 79694
rect 153442 79648 153516 79676
rect 153292 79620 153344 79626
rect 153292 79562 153344 79568
rect 153304 77654 153332 79562
rect 153292 77648 153344 77654
rect 153292 77590 153344 77596
rect 153212 76078 153332 76106
rect 153488 76090 153516 79648
rect 153568 79630 153620 79636
rect 153304 75886 153332 76078
rect 153476 76084 153528 76090
rect 153476 76026 153528 76032
rect 153580 75970 153608 79630
rect 153384 75948 153436 75954
rect 153384 75890 153436 75896
rect 153488 75942 153608 75970
rect 153292 75880 153344 75886
rect 153292 75822 153344 75828
rect 153200 75268 153252 75274
rect 153200 75210 153252 75216
rect 153108 73908 153160 73914
rect 153108 73850 153160 73856
rect 152740 72548 152792 72554
rect 152740 72490 152792 72496
rect 152556 71052 152608 71058
rect 152556 70994 152608 71000
rect 152464 67176 152516 67182
rect 152464 67118 152516 67124
rect 152372 64320 152424 64326
rect 152372 64262 152424 64268
rect 152280 26988 152332 26994
rect 152280 26930 152332 26936
rect 152188 25832 152240 25838
rect 152188 25774 152240 25780
rect 152096 21684 152148 21690
rect 152096 21626 152148 21632
rect 152004 13456 152056 13462
rect 152004 13398 152056 13404
rect 151912 13388 151964 13394
rect 151912 13330 151964 13336
rect 151820 9172 151872 9178
rect 151820 9114 151872 9120
rect 151544 4140 151596 4146
rect 151544 4082 151596 4088
rect 150900 4004 150952 4010
rect 150900 3946 150952 3952
rect 151820 3868 151872 3874
rect 151820 3810 151872 3816
rect 150808 3392 150860 3398
rect 150808 3334 150860 3340
rect 151832 480 151860 3810
rect 152568 3806 152596 70994
rect 153212 70394 153240 75210
rect 153212 70366 153332 70394
rect 153304 5098 153332 70366
rect 153396 13326 153424 75890
rect 153488 23254 153516 75942
rect 153568 75880 153620 75886
rect 153568 75822 153620 75828
rect 153580 31210 153608 75822
rect 153672 65618 153700 79698
rect 153936 79688 153988 79694
rect 153936 79630 153988 79636
rect 153844 79552 153896 79558
rect 153844 79494 153896 79500
rect 153752 79348 153804 79354
rect 153752 79290 153804 79296
rect 153764 68474 153792 79290
rect 153856 77042 153884 79494
rect 153948 79354 153976 79630
rect 153936 79348 153988 79354
rect 153936 79290 153988 79296
rect 154040 78674 154068 79750
rect 154120 79688 154172 79694
rect 154270 79676 154298 80036
rect 154362 79744 154390 80036
rect 154454 79971 154482 80036
rect 154440 79962 154496 79971
rect 154440 79897 154496 79906
rect 154546 79778 154574 80036
rect 154638 79966 154666 80036
rect 154626 79960 154678 79966
rect 154626 79902 154678 79908
rect 154730 79898 154758 80036
rect 154718 79892 154770 79898
rect 154718 79834 154770 79840
rect 154500 79750 154574 79778
rect 154670 79792 154726 79801
rect 154362 79716 154436 79744
rect 154270 79648 154344 79676
rect 154120 79630 154172 79636
rect 153948 78646 154068 78674
rect 153844 77036 153896 77042
rect 153844 76978 153896 76984
rect 153948 75274 153976 78646
rect 154132 75954 154160 79630
rect 154212 79552 154264 79558
rect 154212 79494 154264 79500
rect 154224 78713 154252 79494
rect 154210 78704 154266 78713
rect 154210 78639 154266 78648
rect 154212 78260 154264 78266
rect 154212 78202 154264 78208
rect 154224 77330 154252 78202
rect 154316 78062 154344 79648
rect 154304 78056 154356 78062
rect 154304 77998 154356 78004
rect 154224 77302 154344 77330
rect 154212 77240 154264 77246
rect 154212 77182 154264 77188
rect 154120 75948 154172 75954
rect 154120 75890 154172 75896
rect 153936 75268 153988 75274
rect 153936 75210 153988 75216
rect 153752 68468 153804 68474
rect 153752 68410 153804 68416
rect 153660 65612 153712 65618
rect 153660 65554 153712 65560
rect 154224 64874 154252 77182
rect 154316 70394 154344 77302
rect 154408 75993 154436 79716
rect 154394 75984 154450 75993
rect 154394 75919 154450 75928
rect 154500 75857 154528 79750
rect 154670 79727 154726 79736
rect 154822 79744 154850 80036
rect 154914 79937 154942 80036
rect 155006 79966 155034 80036
rect 155098 79971 155126 80036
rect 154994 79960 155046 79966
rect 154900 79928 154956 79937
rect 154994 79902 155046 79908
rect 155084 79962 155140 79971
rect 155190 79966 155218 80036
rect 155282 79966 155310 80036
rect 155084 79897 155140 79906
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 154900 79863 154956 79872
rect 154948 79824 155000 79830
rect 155374 79812 155402 80036
rect 155466 79898 155494 80036
rect 155558 79971 155586 80036
rect 155544 79962 155600 79971
rect 155454 79892 155506 79898
rect 155544 79897 155600 79906
rect 155454 79834 155506 79840
rect 154948 79766 155000 79772
rect 155038 79792 155094 79801
rect 154580 79688 154632 79694
rect 154580 79630 154632 79636
rect 154592 76226 154620 79630
rect 154684 78266 154712 79727
rect 154822 79716 154896 79744
rect 154764 79620 154816 79626
rect 154764 79562 154816 79568
rect 154672 78260 154724 78266
rect 154672 78202 154724 78208
rect 154580 76220 154632 76226
rect 154580 76162 154632 76168
rect 154672 76152 154724 76158
rect 154672 76094 154724 76100
rect 154580 75948 154632 75954
rect 154580 75890 154632 75896
rect 154486 75848 154542 75857
rect 154486 75783 154542 75792
rect 154316 70366 154528 70394
rect 154132 64846 154252 64874
rect 154132 31278 154160 64846
rect 154120 31272 154172 31278
rect 154120 31214 154172 31220
rect 153568 31204 153620 31210
rect 153568 31146 153620 31152
rect 153476 23248 153528 23254
rect 153476 23190 153528 23196
rect 153384 13320 153436 13326
rect 153384 13262 153436 13268
rect 154500 10538 154528 70366
rect 154592 14618 154620 75890
rect 154684 14754 154712 76094
rect 154776 75818 154804 79562
rect 154868 79354 154896 79716
rect 154856 79348 154908 79354
rect 154856 79290 154908 79296
rect 154960 76548 154988 79766
rect 155038 79727 155094 79736
rect 155144 79784 155402 79812
rect 155052 78946 155080 79727
rect 155144 79490 155172 79784
rect 155650 79778 155678 80036
rect 155742 79937 155770 80036
rect 155728 79928 155784 79937
rect 155834 79898 155862 80036
rect 155926 79898 155954 80036
rect 156018 79966 156046 80036
rect 156006 79960 156058 79966
rect 156110 79937 156138 80036
rect 156006 79902 156058 79908
rect 156096 79928 156152 79937
rect 155728 79863 155784 79872
rect 155822 79892 155874 79898
rect 155822 79834 155874 79840
rect 155914 79892 155966 79898
rect 156202 79898 156230 80036
rect 156294 79966 156322 80036
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156096 79863 156152 79872
rect 156190 79892 156242 79898
rect 155914 79834 155966 79840
rect 156190 79834 156242 79840
rect 156006 79824 156058 79830
rect 155866 79792 155922 79801
rect 155650 79750 155724 79778
rect 155224 79688 155276 79694
rect 155224 79630 155276 79636
rect 155316 79688 155368 79694
rect 155316 79630 155368 79636
rect 155408 79688 155460 79694
rect 155696 79665 155724 79750
rect 155866 79727 155922 79736
rect 155972 79772 156006 79778
rect 156386 79801 156414 80036
rect 156478 79966 156506 80036
rect 156466 79960 156518 79966
rect 156466 79902 156518 79908
rect 156570 79898 156598 80036
rect 156662 79937 156690 80036
rect 156648 79928 156704 79937
rect 156558 79892 156610 79898
rect 156648 79863 156704 79872
rect 156558 79834 156610 79840
rect 156754 79812 156782 80036
rect 156846 79830 156874 80036
rect 156938 79830 156966 80036
rect 157030 79898 157058 80036
rect 157122 79937 157150 80036
rect 157214 79966 157242 80036
rect 157306 79971 157334 80036
rect 157202 79960 157254 79966
rect 157108 79928 157164 79937
rect 157018 79892 157070 79898
rect 157202 79902 157254 79908
rect 157292 79962 157348 79971
rect 157292 79897 157348 79906
rect 157398 79898 157426 80036
rect 157108 79863 157164 79872
rect 157386 79892 157438 79898
rect 157018 79834 157070 79840
rect 157386 79834 157438 79840
rect 155972 79766 156058 79772
rect 156372 79792 156428 79801
rect 155972 79750 156046 79766
rect 155408 79630 155460 79636
rect 155682 79656 155738 79665
rect 155132 79484 155184 79490
rect 155132 79426 155184 79432
rect 155132 79348 155184 79354
rect 155132 79290 155184 79296
rect 155040 78940 155092 78946
rect 155040 78882 155092 78888
rect 155144 78198 155172 79290
rect 155132 78192 155184 78198
rect 155038 78160 155094 78169
rect 155132 78134 155184 78140
rect 155038 78095 155094 78104
rect 154868 76520 154988 76548
rect 154764 75812 154816 75818
rect 154764 75754 154816 75760
rect 154764 75540 154816 75546
rect 154764 75482 154816 75488
rect 154672 14748 154724 14754
rect 154672 14690 154724 14696
rect 154776 14686 154804 75482
rect 154868 16182 154896 76520
rect 155052 75914 155080 78095
rect 155132 76220 155184 76226
rect 155132 76162 155184 76168
rect 154960 75886 155080 75914
rect 154960 23186 154988 75886
rect 155040 75812 155092 75818
rect 155040 75754 155092 75760
rect 155052 24410 155080 75754
rect 155144 63034 155172 76162
rect 155236 76158 155264 79630
rect 155224 76152 155276 76158
rect 155224 76094 155276 76100
rect 155222 75984 155278 75993
rect 155222 75919 155278 75928
rect 155236 65550 155264 75919
rect 155328 70038 155356 79630
rect 155420 75546 155448 79630
rect 155682 79591 155738 79600
rect 155776 79484 155828 79490
rect 155776 79426 155828 79432
rect 155500 78940 155552 78946
rect 155500 78882 155552 78888
rect 155512 75954 155540 78882
rect 155788 76294 155816 79426
rect 155776 76288 155828 76294
rect 155880 76265 155908 79727
rect 155776 76230 155828 76236
rect 155866 76256 155922 76265
rect 155866 76191 155922 76200
rect 155868 76084 155920 76090
rect 155868 76026 155920 76032
rect 155500 75948 155552 75954
rect 155500 75890 155552 75896
rect 155408 75540 155460 75546
rect 155408 75482 155460 75488
rect 155880 72486 155908 76026
rect 155972 75886 156000 79750
rect 156708 79784 156782 79812
rect 156834 79824 156886 79830
rect 156372 79727 156428 79736
rect 156512 79756 156564 79762
rect 156512 79698 156564 79704
rect 156604 79756 156656 79762
rect 156604 79698 156656 79704
rect 156144 79688 156196 79694
rect 156050 79656 156106 79665
rect 156144 79630 156196 79636
rect 156050 79591 156106 79600
rect 156064 76362 156092 79591
rect 156156 77994 156184 79630
rect 156236 79620 156288 79626
rect 156236 79562 156288 79568
rect 156144 77988 156196 77994
rect 156144 77930 156196 77936
rect 156144 77852 156196 77858
rect 156144 77794 156196 77800
rect 156156 77314 156184 77794
rect 156144 77308 156196 77314
rect 156144 77250 156196 77256
rect 156052 76356 156104 76362
rect 156052 76298 156104 76304
rect 156248 76242 156276 79562
rect 156328 79552 156380 79558
rect 156328 79494 156380 79500
rect 156064 76214 156276 76242
rect 155960 75880 156012 75886
rect 155960 75822 156012 75828
rect 155960 75404 156012 75410
rect 155960 75346 156012 75352
rect 155868 72480 155920 72486
rect 155868 72422 155920 72428
rect 155316 70032 155368 70038
rect 155316 69974 155368 69980
rect 155224 65544 155276 65550
rect 155224 65486 155276 65492
rect 155132 63028 155184 63034
rect 155132 62970 155184 62976
rect 155040 24404 155092 24410
rect 155040 24346 155092 24352
rect 154948 23180 155000 23186
rect 154948 23122 155000 23128
rect 154856 16176 154908 16182
rect 154856 16118 154908 16124
rect 154764 14680 154816 14686
rect 154764 14622 154816 14628
rect 154580 14612 154632 14618
rect 154580 14554 154632 14560
rect 154488 10532 154540 10538
rect 154488 10474 154540 10480
rect 155972 7818 156000 75346
rect 156064 10470 156092 76214
rect 156236 76084 156288 76090
rect 156236 76026 156288 76032
rect 156142 75984 156198 75993
rect 156142 75919 156198 75928
rect 156052 10464 156104 10470
rect 156052 10406 156104 10412
rect 156156 10402 156184 75919
rect 156248 16046 156276 76026
rect 156340 16114 156368 79494
rect 156420 79484 156472 79490
rect 156420 79426 156472 79432
rect 156432 77897 156460 79426
rect 156418 77888 156474 77897
rect 156418 77823 156474 77832
rect 156420 76356 156472 76362
rect 156420 76298 156472 76304
rect 156432 32774 156460 76298
rect 156524 76090 156552 79698
rect 156512 76084 156564 76090
rect 156512 76026 156564 76032
rect 156616 75970 156644 79698
rect 156524 75942 156644 75970
rect 156524 58682 156552 75942
rect 156604 75880 156656 75886
rect 156604 75822 156656 75828
rect 156616 69970 156644 75822
rect 156708 75410 156736 79784
rect 156834 79766 156886 79772
rect 156926 79824 156978 79830
rect 156926 79766 156978 79772
rect 157156 79824 157208 79830
rect 157156 79766 157208 79772
rect 156880 79688 156932 79694
rect 156786 79656 156842 79665
rect 156880 79630 156932 79636
rect 156786 79591 156842 79600
rect 156800 75818 156828 79591
rect 156788 75812 156840 75818
rect 156788 75754 156840 75760
rect 156892 75449 156920 79630
rect 157064 79620 157116 79626
rect 157064 79562 157116 79568
rect 156972 79416 157024 79422
rect 156972 79358 157024 79364
rect 156878 75440 156934 75449
rect 156696 75404 156748 75410
rect 156878 75375 156934 75384
rect 156696 75346 156748 75352
rect 156604 69964 156656 69970
rect 156604 69906 156656 69912
rect 156512 58676 156564 58682
rect 156512 58618 156564 58624
rect 156420 32768 156472 32774
rect 156420 32710 156472 32716
rect 156984 31142 157012 79358
rect 157076 77489 157104 79562
rect 157168 78305 157196 79766
rect 157490 79676 157518 80036
rect 157582 79744 157610 80036
rect 157674 79898 157702 80036
rect 157766 79966 157794 80036
rect 157858 79966 157886 80036
rect 157754 79960 157806 79966
rect 157754 79902 157806 79908
rect 157846 79960 157898 79966
rect 157846 79902 157898 79908
rect 157662 79892 157714 79898
rect 157662 79834 157714 79840
rect 157950 79778 157978 80036
rect 158042 79966 158070 80036
rect 158030 79960 158082 79966
rect 158030 79902 158082 79908
rect 157950 79750 158024 79778
rect 157582 79716 157656 79744
rect 157444 79648 157518 79676
rect 157340 79620 157392 79626
rect 157340 79562 157392 79568
rect 157248 79008 157300 79014
rect 157248 78950 157300 78956
rect 157260 78849 157288 78950
rect 157246 78840 157302 78849
rect 157246 78775 157302 78784
rect 157154 78296 157210 78305
rect 157154 78231 157210 78240
rect 157062 77480 157118 77489
rect 157062 77415 157118 77424
rect 157064 77308 157116 77314
rect 157064 77250 157116 77256
rect 157076 68542 157104 77250
rect 157352 76684 157380 79562
rect 157260 76656 157380 76684
rect 157260 75954 157288 76656
rect 157444 76616 157472 79648
rect 157524 79552 157576 79558
rect 157524 79494 157576 79500
rect 157352 76588 157472 76616
rect 157248 75948 157300 75954
rect 157248 75890 157300 75896
rect 157064 68536 157116 68542
rect 157064 68478 157116 68484
rect 156972 31136 157024 31142
rect 156972 31078 157024 31084
rect 156328 16108 156380 16114
rect 156328 16050 156380 16056
rect 156236 16040 156288 16046
rect 156236 15982 156288 15988
rect 156144 10396 156196 10402
rect 156144 10338 156196 10344
rect 155960 7812 156012 7818
rect 155960 7754 156012 7760
rect 157352 6526 157380 76588
rect 157536 75914 157564 79494
rect 157628 79422 157656 79716
rect 157708 79620 157760 79626
rect 157892 79620 157944 79626
rect 157760 79580 157840 79608
rect 157708 79562 157760 79568
rect 157616 79416 157668 79422
rect 157616 79358 157668 79364
rect 157708 78940 157760 78946
rect 157708 78882 157760 78888
rect 157616 78804 157668 78810
rect 157616 78746 157668 78752
rect 157444 75886 157564 75914
rect 157444 11898 157472 75886
rect 157524 75268 157576 75274
rect 157524 75210 157576 75216
rect 157432 11892 157484 11898
rect 157432 11834 157484 11840
rect 157536 11830 157564 75210
rect 157628 13258 157656 78746
rect 157720 17610 157748 78882
rect 157812 78112 157840 79580
rect 157892 79562 157944 79568
rect 157904 78674 157932 79562
rect 157996 78946 158024 79750
rect 158134 79744 158162 80036
rect 158226 79966 158254 80036
rect 158318 79966 158346 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158306 79960 158358 79966
rect 158410 79937 158438 80036
rect 158502 79966 158530 80036
rect 158490 79960 158542 79966
rect 158306 79902 158358 79908
rect 158396 79928 158452 79937
rect 158594 79937 158622 80036
rect 158490 79902 158542 79908
rect 158580 79928 158636 79937
rect 158396 79863 158452 79872
rect 158580 79863 158636 79872
rect 158444 79756 158496 79762
rect 158134 79716 158208 79744
rect 158180 79676 158208 79716
rect 158686 79744 158714 80036
rect 158778 79966 158806 80036
rect 158870 79966 158898 80036
rect 158962 79971 158990 80036
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158858 79960 158910 79966
rect 158858 79902 158910 79908
rect 158948 79962 159004 79971
rect 159054 79966 159082 80036
rect 158948 79897 159004 79906
rect 159042 79960 159094 79966
rect 159042 79902 159094 79908
rect 158858 79824 158910 79830
rect 159146 79778 159174 80036
rect 159238 79966 159266 80036
rect 159330 79966 159358 80036
rect 159226 79960 159278 79966
rect 159226 79902 159278 79908
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 159422 79898 159450 80036
rect 159514 79966 159542 80036
rect 159606 79966 159634 80036
rect 159502 79960 159554 79966
rect 159502 79902 159554 79908
rect 159594 79960 159646 79966
rect 159594 79902 159646 79908
rect 159698 79898 159726 80036
rect 159790 79971 159818 80036
rect 159776 79962 159832 79971
rect 159410 79892 159462 79898
rect 159410 79834 159462 79840
rect 159686 79892 159738 79898
rect 159776 79897 159832 79906
rect 159686 79834 159738 79840
rect 158858 79766 158910 79772
rect 158444 79698 158496 79704
rect 158640 79716 158714 79744
rect 158180 79648 158392 79676
rect 158076 79620 158128 79626
rect 158076 79562 158128 79568
rect 157984 78940 158036 78946
rect 157984 78882 158036 78888
rect 158088 78810 158116 79562
rect 158168 79552 158220 79558
rect 158168 79494 158220 79500
rect 158076 78804 158128 78810
rect 158076 78746 158128 78752
rect 157892 78668 157944 78674
rect 157892 78610 157944 78616
rect 158076 78668 158128 78674
rect 158076 78610 158128 78616
rect 157812 78084 157932 78112
rect 157800 75200 157852 75206
rect 157800 75142 157852 75148
rect 157708 17604 157760 17610
rect 157708 17546 157760 17552
rect 157812 17542 157840 75142
rect 157904 61470 157932 78084
rect 158088 75274 158116 78610
rect 158076 75268 158128 75274
rect 158076 75210 158128 75216
rect 158180 75206 158208 79494
rect 158364 77722 158392 79648
rect 158456 78033 158484 79698
rect 158536 79688 158588 79694
rect 158536 79630 158588 79636
rect 158548 78169 158576 79630
rect 158534 78160 158590 78169
rect 158534 78095 158590 78104
rect 158442 78024 158498 78033
rect 158442 77959 158498 77968
rect 158640 77858 158668 79716
rect 158870 79676 158898 79766
rect 158732 79648 158898 79676
rect 159008 79750 159174 79778
rect 159732 79756 159784 79762
rect 158628 77852 158680 77858
rect 158628 77794 158680 77800
rect 158352 77716 158404 77722
rect 158352 77658 158404 77664
rect 158260 77444 158312 77450
rect 158260 77386 158312 77392
rect 158272 77194 158300 77386
rect 158272 77166 158392 77194
rect 158260 75948 158312 75954
rect 158260 75890 158312 75896
rect 158168 75200 158220 75206
rect 158168 75142 158220 75148
rect 158272 70394 158300 75890
rect 158364 71058 158392 77166
rect 158732 76566 158760 79648
rect 158904 79552 158956 79558
rect 158904 79494 158956 79500
rect 158810 78568 158866 78577
rect 158810 78503 158866 78512
rect 158720 76560 158772 76566
rect 158720 76502 158772 76508
rect 158720 76356 158772 76362
rect 158720 76298 158772 76304
rect 158352 71052 158404 71058
rect 158352 70994 158404 71000
rect 158088 70366 158300 70394
rect 158088 64874 158116 70366
rect 157996 64846 158116 64874
rect 157996 62966 158024 64846
rect 157984 62960 158036 62966
rect 157984 62902 158036 62908
rect 157892 61464 157944 61470
rect 157892 61406 157944 61412
rect 157800 17536 157852 17542
rect 157800 17478 157852 17484
rect 157616 13252 157668 13258
rect 157616 13194 157668 13200
rect 157524 11824 157576 11830
rect 157524 11766 157576 11772
rect 157340 6520 157392 6526
rect 157340 6462 157392 6468
rect 158732 6390 158760 76298
rect 158824 13190 158852 78503
rect 158916 14550 158944 79494
rect 159008 75682 159036 79750
rect 159732 79698 159784 79704
rect 159088 79688 159140 79694
rect 159088 79630 159140 79636
rect 159364 79688 159416 79694
rect 159364 79630 159416 79636
rect 158996 75676 159048 75682
rect 158996 75618 159048 75624
rect 159100 60042 159128 79630
rect 159180 79620 159232 79626
rect 159180 79562 159232 79568
rect 159272 79620 159324 79626
rect 159272 79562 159324 79568
rect 159192 78878 159220 79562
rect 159180 78872 159232 78878
rect 159180 78814 159232 78820
rect 159180 78736 159232 78742
rect 159180 78678 159232 78684
rect 159192 78033 159220 78678
rect 159178 78024 159234 78033
rect 159178 77959 159234 77968
rect 159284 77790 159312 79562
rect 159376 79506 159404 79630
rect 159376 79478 159496 79506
rect 159364 78940 159416 78946
rect 159364 78882 159416 78888
rect 159272 77784 159324 77790
rect 159272 77726 159324 77732
rect 159376 76650 159404 78882
rect 159192 76622 159404 76650
rect 159192 67114 159220 76622
rect 159468 76566 159496 79478
rect 159640 79348 159692 79354
rect 159640 79290 159692 79296
rect 159652 78130 159680 79290
rect 159744 78713 159772 79698
rect 159882 79642 159910 80036
rect 159974 79898 160002 80036
rect 160066 79971 160094 80036
rect 160052 79962 160108 79971
rect 159962 79892 160014 79898
rect 160052 79897 160108 79906
rect 160158 79898 160186 80036
rect 159962 79834 160014 79840
rect 160146 79892 160198 79898
rect 160146 79834 160198 79840
rect 160250 79744 160278 80036
rect 160342 79966 160370 80036
rect 160434 79966 160462 80036
rect 160526 79971 160554 80036
rect 160330 79960 160382 79966
rect 160330 79902 160382 79908
rect 160422 79960 160474 79966
rect 160422 79902 160474 79908
rect 160512 79962 160568 79971
rect 160512 79897 160568 79906
rect 160618 79898 160646 80036
rect 160710 79966 160738 80036
rect 160698 79960 160750 79966
rect 160698 79902 160750 79908
rect 160606 79892 160658 79898
rect 160606 79834 160658 79840
rect 160468 79824 160520 79830
rect 160468 79766 160520 79772
rect 160204 79716 160278 79744
rect 160376 79756 160428 79762
rect 159836 79614 159910 79642
rect 160008 79688 160060 79694
rect 160008 79630 160060 79636
rect 159730 78704 159786 78713
rect 159730 78639 159786 78648
rect 159640 78124 159692 78130
rect 159640 78066 159692 78072
rect 159836 77294 159864 79614
rect 159916 79416 159968 79422
rect 159916 79358 159968 79364
rect 159928 77654 159956 79358
rect 159916 77648 159968 77654
rect 159916 77590 159968 77596
rect 159744 77266 159864 77294
rect 159272 76560 159324 76566
rect 159272 76502 159324 76508
rect 159456 76560 159508 76566
rect 159456 76502 159508 76508
rect 159284 68406 159312 76502
rect 159744 76362 159772 77266
rect 160020 76650 160048 79630
rect 160204 78928 160232 79716
rect 160376 79698 160428 79704
rect 160284 79620 160336 79626
rect 160284 79562 160336 79568
rect 160296 78946 160324 79562
rect 159928 76622 160048 76650
rect 160112 78900 160232 78928
rect 160284 78940 160336 78946
rect 159732 76356 159784 76362
rect 159732 76298 159784 76304
rect 159640 76288 159692 76294
rect 159640 76230 159692 76236
rect 159652 70394 159680 76230
rect 159928 75614 159956 76622
rect 160008 76560 160060 76566
rect 160008 76502 160060 76508
rect 159916 75608 159968 75614
rect 159916 75550 159968 75556
rect 159652 70366 159772 70394
rect 159272 68400 159324 68406
rect 159272 68342 159324 68348
rect 159180 67108 159232 67114
rect 159180 67050 159232 67056
rect 159088 60036 159140 60042
rect 159088 59978 159140 59984
rect 159744 35222 159772 70366
rect 159732 35216 159784 35222
rect 159732 35158 159784 35164
rect 160020 32706 160048 76502
rect 160008 32700 160060 32706
rect 160008 32642 160060 32648
rect 158904 14544 158956 14550
rect 158904 14486 158956 14492
rect 158812 13184 158864 13190
rect 158812 13126 158864 13132
rect 160112 7750 160140 78900
rect 160284 78882 160336 78888
rect 160192 78804 160244 78810
rect 160192 78746 160244 78752
rect 160204 76566 160232 78746
rect 160282 78704 160338 78713
rect 160282 78639 160338 78648
rect 160192 76560 160244 76566
rect 160192 76502 160244 76508
rect 160192 75200 160244 75206
rect 160192 75142 160244 75148
rect 160204 13122 160232 75142
rect 160296 17406 160324 78639
rect 160388 77586 160416 79698
rect 160376 77580 160428 77586
rect 160376 77522 160428 77528
rect 160376 75268 160428 75274
rect 160376 75210 160428 75216
rect 160388 18834 160416 75210
rect 160480 18902 160508 79766
rect 160560 79688 160612 79694
rect 160802 79676 160830 80036
rect 160894 79971 160922 80036
rect 160880 79962 160936 79971
rect 160880 79897 160936 79906
rect 160986 79898 161014 80036
rect 161078 79966 161106 80036
rect 161170 79966 161198 80036
rect 161262 79966 161290 80036
rect 161354 79971 161382 80036
rect 161066 79960 161118 79966
rect 161066 79902 161118 79908
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161250 79960 161302 79966
rect 161250 79902 161302 79908
rect 161340 79962 161396 79971
rect 160974 79892 161026 79898
rect 161340 79897 161396 79906
rect 160974 79834 161026 79840
rect 161446 79830 161474 80036
rect 161538 79971 161566 80036
rect 161524 79962 161580 79971
rect 161524 79897 161580 79906
rect 161630 79898 161658 80036
rect 161618 79892 161670 79898
rect 161618 79834 161670 79840
rect 161434 79824 161486 79830
rect 161294 79792 161350 79801
rect 161020 79756 161072 79762
rect 161020 79698 161072 79704
rect 161112 79756 161164 79762
rect 161722 79778 161750 80036
rect 161814 79966 161842 80036
rect 161906 79966 161934 80036
rect 161802 79960 161854 79966
rect 161802 79902 161854 79908
rect 161894 79960 161946 79966
rect 161998 79937 162026 80036
rect 162090 79966 162118 80036
rect 162078 79960 162130 79966
rect 161894 79902 161946 79908
rect 161984 79928 162040 79937
rect 162078 79902 162130 79908
rect 161984 79863 162040 79872
rect 161434 79766 161486 79772
rect 161294 79727 161350 79736
rect 161572 79756 161624 79762
rect 161112 79698 161164 79704
rect 160560 79630 160612 79636
rect 160756 79648 160830 79676
rect 160926 79656 160982 79665
rect 160572 79082 160600 79630
rect 160652 79620 160704 79626
rect 160652 79562 160704 79568
rect 160560 79076 160612 79082
rect 160560 79018 160612 79024
rect 160560 78668 160612 78674
rect 160560 78610 160612 78616
rect 160572 20058 160600 78610
rect 160664 77994 160692 79562
rect 160756 78554 160784 79648
rect 160926 79591 160982 79600
rect 160836 79552 160888 79558
rect 160836 79494 160888 79500
rect 160848 78674 160876 79494
rect 160940 78810 160968 79591
rect 160928 78804 160980 78810
rect 160928 78746 160980 78752
rect 161032 78713 161060 79698
rect 161018 78704 161074 78713
rect 160836 78668 160888 78674
rect 160836 78610 160888 78616
rect 160928 78668 160980 78674
rect 161018 78639 161074 78648
rect 160928 78610 160980 78616
rect 160756 78526 160876 78554
rect 160744 78260 160796 78266
rect 160744 78202 160796 78208
rect 160652 77988 160704 77994
rect 160652 77930 160704 77936
rect 160652 77580 160704 77586
rect 160652 77522 160704 77528
rect 160664 21622 160692 77522
rect 160756 75274 160784 78202
rect 160744 75268 160796 75274
rect 160744 75210 160796 75216
rect 160848 75206 160876 78526
rect 160940 78470 160968 78610
rect 160928 78464 160980 78470
rect 160928 78406 160980 78412
rect 161124 78334 161152 79698
rect 161204 79688 161256 79694
rect 161204 79630 161256 79636
rect 161216 78577 161244 79630
rect 161308 79626 161336 79727
rect 161572 79698 161624 79704
rect 161676 79750 161750 79778
rect 161940 79824 161992 79830
rect 161940 79766 161992 79772
rect 161848 79756 161900 79762
rect 161480 79688 161532 79694
rect 161386 79656 161442 79665
rect 161296 79620 161348 79626
rect 161480 79630 161532 79636
rect 161386 79591 161442 79600
rect 161296 79562 161348 79568
rect 161296 79076 161348 79082
rect 161296 79018 161348 79024
rect 161202 78568 161258 78577
rect 161202 78503 161258 78512
rect 161204 78464 161256 78470
rect 161204 78406 161256 78412
rect 160928 78328 160980 78334
rect 160928 78270 160980 78276
rect 161112 78328 161164 78334
rect 161112 78270 161164 78276
rect 160836 75200 160888 75206
rect 160836 75142 160888 75148
rect 160940 70394 160968 78270
rect 161020 78192 161072 78198
rect 161020 78134 161072 78140
rect 161032 73846 161060 78134
rect 161216 78033 161244 78406
rect 161308 78266 161336 79018
rect 161296 78260 161348 78266
rect 161296 78202 161348 78208
rect 161202 78024 161258 78033
rect 161202 77959 161258 77968
rect 161400 75914 161428 79591
rect 161492 78441 161520 79630
rect 161584 78810 161612 79698
rect 161676 79558 161704 79750
rect 161848 79698 161900 79704
rect 161756 79688 161808 79694
rect 161860 79665 161888 79698
rect 161756 79630 161808 79636
rect 161846 79656 161902 79665
rect 161664 79552 161716 79558
rect 161664 79494 161716 79500
rect 161664 78940 161716 78946
rect 161664 78882 161716 78888
rect 161572 78804 161624 78810
rect 161572 78746 161624 78752
rect 161570 78704 161626 78713
rect 161570 78639 161626 78648
rect 161478 78432 161534 78441
rect 161478 78367 161534 78376
rect 161400 75886 161520 75914
rect 161020 73840 161072 73846
rect 161020 73782 161072 73788
rect 160848 70366 160968 70394
rect 160848 67250 160876 70366
rect 160836 67244 160888 67250
rect 160836 67186 160888 67192
rect 160652 21616 160704 21622
rect 160652 21558 160704 21564
rect 160560 20052 160612 20058
rect 160560 19994 160612 20000
rect 160558 19952 160614 19961
rect 160558 19887 160614 19896
rect 160468 18896 160520 18902
rect 160468 18838 160520 18844
rect 160376 18828 160428 18834
rect 160376 18770 160428 18776
rect 160284 17400 160336 17406
rect 160284 17342 160336 17348
rect 160192 13116 160244 13122
rect 160192 13058 160244 13064
rect 160100 7744 160152 7750
rect 160100 7686 160152 7692
rect 160572 6914 160600 19887
rect 160112 6886 160600 6914
rect 158720 6384 158772 6390
rect 158720 6326 158772 6332
rect 156604 6248 156656 6254
rect 156604 6190 156656 6196
rect 153292 5092 153344 5098
rect 153292 5034 153344 5040
rect 152556 3800 152608 3806
rect 152556 3742 152608 3748
rect 154212 3732 154264 3738
rect 154212 3674 154264 3680
rect 153016 3324 153068 3330
rect 153016 3266 153068 3272
rect 153028 480 153056 3266
rect 154224 480 154252 3674
rect 155408 3664 155460 3670
rect 155408 3606 155460 3612
rect 155420 480 155448 3606
rect 156616 480 156644 6190
rect 157800 4888 157852 4894
rect 157800 4830 157852 4836
rect 158902 4856 158958 4865
rect 157812 480 157840 4830
rect 158902 4791 158958 4800
rect 158916 480 158944 4791
rect 160112 480 160140 6886
rect 161492 6322 161520 75886
rect 161584 75274 161612 78639
rect 161572 75268 161624 75274
rect 161572 75210 161624 75216
rect 161572 75132 161624 75138
rect 161572 75074 161624 75080
rect 161584 7682 161612 75074
rect 161676 9110 161704 78882
rect 161768 19990 161796 79630
rect 161846 79591 161902 79600
rect 161848 79484 161900 79490
rect 161848 79426 161900 79432
rect 161860 79150 161888 79426
rect 161952 79354 161980 79766
rect 162032 79756 162084 79762
rect 162182 79744 162210 80036
rect 162274 79898 162302 80036
rect 162366 79898 162394 80036
rect 162458 79898 162486 80036
rect 162262 79892 162314 79898
rect 162262 79834 162314 79840
rect 162354 79892 162406 79898
rect 162354 79834 162406 79840
rect 162446 79892 162498 79898
rect 162446 79834 162498 79840
rect 162398 79792 162454 79801
rect 162182 79716 162256 79744
rect 162398 79727 162454 79736
rect 162550 79744 162578 80036
rect 162642 79937 162670 80036
rect 162628 79928 162684 79937
rect 162628 79863 162684 79872
rect 162734 79801 162762 80036
rect 162720 79792 162776 79801
rect 162032 79698 162084 79704
rect 161940 79348 161992 79354
rect 161940 79290 161992 79296
rect 161848 79144 161900 79150
rect 161848 79086 161900 79092
rect 161940 78804 161992 78810
rect 161940 78746 161992 78752
rect 161848 78736 161900 78742
rect 161848 78678 161900 78684
rect 161860 21554 161888 78678
rect 161952 32638 161980 78746
rect 162044 77294 162072 79698
rect 162124 79620 162176 79626
rect 162124 79562 162176 79568
rect 162136 78742 162164 79562
rect 162228 78946 162256 79716
rect 162308 79688 162360 79694
rect 162308 79630 162360 79636
rect 162412 79642 162440 79727
rect 162550 79716 162624 79744
rect 162826 79778 162854 80036
rect 162918 79898 162946 80036
rect 163010 79971 163038 80036
rect 162996 79962 163052 79971
rect 162906 79892 162958 79898
rect 162996 79897 163052 79906
rect 162906 79834 162958 79840
rect 162950 79792 163006 79801
rect 162826 79750 162900 79778
rect 162720 79727 162776 79736
rect 162216 78940 162268 78946
rect 162216 78882 162268 78888
rect 162216 78804 162268 78810
rect 162216 78746 162268 78752
rect 162124 78736 162176 78742
rect 162124 78678 162176 78684
rect 162122 78432 162178 78441
rect 162122 78367 162178 78376
rect 162136 78130 162164 78367
rect 162124 78124 162176 78130
rect 162124 78066 162176 78072
rect 162228 77382 162256 78746
rect 162320 78130 162348 79630
rect 162412 79626 162532 79642
rect 162412 79620 162544 79626
rect 162412 79614 162492 79620
rect 162492 79562 162544 79568
rect 162400 79552 162452 79558
rect 162400 79494 162452 79500
rect 162412 78266 162440 79494
rect 162596 79064 162624 79716
rect 162676 79688 162728 79694
rect 162676 79630 162728 79636
rect 162768 79688 162820 79694
rect 162768 79630 162820 79636
rect 162504 79036 162624 79064
rect 162504 78713 162532 79036
rect 162584 78940 162636 78946
rect 162584 78882 162636 78888
rect 162490 78704 162546 78713
rect 162490 78639 162546 78648
rect 162400 78260 162452 78266
rect 162400 78202 162452 78208
rect 162308 78124 162360 78130
rect 162308 78066 162360 78072
rect 162400 78056 162452 78062
rect 162400 77998 162452 78004
rect 162308 77920 162360 77926
rect 162308 77862 162360 77868
rect 162216 77376 162268 77382
rect 162216 77318 162268 77324
rect 162044 77266 162164 77294
rect 162032 75268 162084 75274
rect 162032 75210 162084 75216
rect 162044 67046 162072 75210
rect 162136 75138 162164 77266
rect 162214 77208 162270 77217
rect 162214 77143 162270 77152
rect 162228 75546 162256 77143
rect 162216 75540 162268 75546
rect 162216 75482 162268 75488
rect 162124 75132 162176 75138
rect 162124 75074 162176 75080
rect 162032 67040 162084 67046
rect 162032 66982 162084 66988
rect 162320 64874 162348 77862
rect 162412 70394 162440 77998
rect 162596 77294 162624 78882
rect 162688 78713 162716 79630
rect 162674 78704 162730 78713
rect 162674 78639 162730 78648
rect 162780 78062 162808 79630
rect 162768 78056 162820 78062
rect 162872 78033 162900 79750
rect 163102 79744 163130 80036
rect 163194 79971 163222 80036
rect 163180 79962 163236 79971
rect 163180 79897 163236 79906
rect 163286 79898 163314 80036
rect 163274 79892 163326 79898
rect 163274 79834 163326 79840
rect 163378 79801 163406 80036
rect 163470 79812 163498 80036
rect 163562 79971 163590 80036
rect 163548 79962 163604 79971
rect 163548 79897 163604 79906
rect 163654 79898 163682 80036
rect 163746 79898 163774 80036
rect 163838 79937 163866 80036
rect 163930 79966 163958 80036
rect 164022 79971 164050 80036
rect 163918 79960 163970 79966
rect 163824 79928 163880 79937
rect 163642 79892 163694 79898
rect 163642 79834 163694 79840
rect 163734 79892 163786 79898
rect 163918 79902 163970 79908
rect 164008 79962 164064 79971
rect 164008 79897 164064 79906
rect 163824 79863 163880 79872
rect 163734 79834 163786 79840
rect 163964 79824 164016 79830
rect 163364 79792 163420 79801
rect 162950 79727 163006 79736
rect 162964 78946 162992 79727
rect 163056 79716 163130 79744
rect 163228 79756 163280 79762
rect 162952 78940 163004 78946
rect 162952 78882 163004 78888
rect 162952 78192 163004 78198
rect 162952 78134 163004 78140
rect 162768 77998 162820 78004
rect 162858 78024 162914 78033
rect 162858 77959 162914 77968
rect 162596 77266 162900 77294
rect 162872 75206 162900 77266
rect 162860 75200 162912 75206
rect 162860 75142 162912 75148
rect 162412 70366 162624 70394
rect 162228 64846 162348 64874
rect 162228 42090 162256 64846
rect 162596 64258 162624 70366
rect 162584 64252 162636 64258
rect 162584 64194 162636 64200
rect 162216 42084 162268 42090
rect 162216 42026 162268 42032
rect 161940 32632 161992 32638
rect 161940 32574 161992 32580
rect 161848 21548 161900 21554
rect 161848 21490 161900 21496
rect 162860 20120 162912 20126
rect 162860 20062 162912 20068
rect 161756 19984 161808 19990
rect 161756 19926 161808 19932
rect 161664 9104 161716 9110
rect 161664 9046 161716 9052
rect 161572 7676 161624 7682
rect 161572 7618 161624 7624
rect 161480 6316 161532 6322
rect 161480 6258 161532 6264
rect 162492 6180 162544 6186
rect 162492 6122 162544 6128
rect 161294 3360 161350 3369
rect 161294 3295 161350 3304
rect 161308 480 161336 3295
rect 162504 480 162532 6122
rect 162872 3482 162900 20062
rect 162964 4962 162992 78134
rect 163056 75274 163084 79716
rect 163470 79784 163590 79812
rect 163562 79778 163590 79784
rect 163870 79792 163926 79801
rect 163562 79750 163636 79778
rect 163364 79727 163420 79736
rect 163608 79744 163636 79750
rect 163780 79756 163832 79762
rect 163608 79716 163728 79744
rect 163228 79698 163280 79704
rect 163136 79552 163188 79558
rect 163136 79494 163188 79500
rect 163148 78470 163176 79494
rect 163240 78713 163268 79698
rect 163320 79688 163372 79694
rect 163320 79630 163372 79636
rect 163412 79688 163464 79694
rect 163412 79630 163464 79636
rect 163226 78704 163282 78713
rect 163226 78639 163282 78648
rect 163136 78464 163188 78470
rect 163136 78406 163188 78412
rect 163228 77920 163280 77926
rect 163228 77862 163280 77868
rect 163134 77616 163190 77625
rect 163134 77551 163190 77560
rect 163044 75268 163096 75274
rect 163044 75210 163096 75216
rect 163044 75132 163096 75138
rect 163044 75074 163096 75080
rect 163056 9042 163084 75074
rect 163148 10334 163176 77551
rect 163240 17338 163268 77862
rect 163332 21486 163360 79630
rect 163424 79558 163452 79630
rect 163412 79552 163464 79558
rect 163412 79494 163464 79500
rect 163412 79348 163464 79354
rect 163412 79290 163464 79296
rect 163424 77382 163452 79290
rect 163504 79144 163556 79150
rect 163504 79086 163556 79092
rect 163516 78849 163544 79086
rect 163700 79064 163728 79716
rect 164114 79812 164142 80036
rect 164206 79966 164234 80036
rect 164194 79960 164246 79966
rect 164298 79937 164326 80036
rect 164194 79902 164246 79908
rect 164284 79928 164340 79937
rect 164284 79863 164340 79872
rect 164114 79784 164188 79812
rect 163964 79766 164016 79772
rect 164160 79778 164188 79784
rect 163870 79727 163926 79736
rect 163780 79698 163832 79704
rect 163608 79036 163728 79064
rect 163502 78840 163558 78849
rect 163502 78775 163558 78784
rect 163608 78198 163636 79036
rect 163596 78192 163648 78198
rect 163596 78134 163648 78140
rect 163594 77752 163650 77761
rect 163594 77687 163650 77696
rect 163412 77376 163464 77382
rect 163412 77318 163464 77324
rect 163412 75268 163464 75274
rect 163412 75210 163464 75216
rect 163424 32570 163452 75210
rect 163504 75200 163556 75206
rect 163504 75142 163556 75148
rect 163516 57322 163544 75142
rect 163608 62898 163636 77687
rect 163792 70394 163820 79698
rect 163884 75138 163912 79727
rect 163976 79642 164004 79766
rect 164160 79750 164280 79778
rect 164148 79688 164200 79694
rect 163976 79614 164096 79642
rect 164252 79665 164280 79750
rect 164390 79676 164418 80036
rect 164482 79744 164510 80036
rect 164574 79971 164602 80036
rect 164560 79962 164616 79971
rect 164560 79897 164616 79906
rect 164666 79744 164694 80036
rect 164758 79812 164786 80036
rect 164850 79966 164878 80036
rect 164942 79966 164970 80036
rect 164838 79960 164890 79966
rect 164838 79902 164890 79908
rect 164930 79960 164982 79966
rect 164930 79902 164982 79908
rect 164758 79784 164832 79812
rect 164482 79716 164556 79744
rect 164666 79716 164740 79744
rect 164148 79630 164200 79636
rect 164238 79656 164294 79665
rect 163964 79552 164016 79558
rect 163964 79494 164016 79500
rect 163976 75478 164004 79494
rect 164068 77926 164096 79614
rect 164056 77920 164108 77926
rect 164056 77862 164108 77868
rect 163964 75472 164016 75478
rect 163964 75414 164016 75420
rect 164160 75313 164188 79630
rect 164390 79648 164464 79676
rect 164238 79591 164294 79600
rect 164332 79552 164384 79558
rect 164332 79494 164384 79500
rect 164240 78940 164292 78946
rect 164240 78882 164292 78888
rect 164146 75304 164202 75313
rect 164146 75239 164202 75248
rect 163872 75132 163924 75138
rect 163872 75074 163924 75080
rect 163792 70366 164004 70394
rect 163596 62892 163648 62898
rect 163596 62834 163648 62840
rect 163504 57316 163556 57322
rect 163504 57258 163556 57264
rect 163412 32564 163464 32570
rect 163412 32506 163464 32512
rect 163320 21480 163372 21486
rect 163320 21422 163372 21428
rect 163228 17332 163280 17338
rect 163228 17274 163280 17280
rect 163136 10328 163188 10334
rect 163136 10270 163188 10276
rect 163044 9036 163096 9042
rect 163044 8978 163096 8984
rect 162952 4956 163004 4962
rect 162952 4898 163004 4904
rect 163976 3738 164004 70366
rect 164252 7614 164280 78882
rect 164344 14482 164372 79494
rect 164436 75914 164464 79648
rect 164528 79608 164556 79716
rect 164712 79626 164740 79716
rect 164700 79620 164752 79626
rect 164528 79580 164648 79608
rect 164516 79484 164568 79490
rect 164516 79426 164568 79432
rect 164528 79286 164556 79426
rect 164516 79280 164568 79286
rect 164516 79222 164568 79228
rect 164516 79008 164568 79014
rect 164516 78950 164568 78956
rect 164528 78742 164556 78950
rect 164516 78736 164568 78742
rect 164516 78678 164568 78684
rect 164436 75886 164556 75914
rect 164424 75404 164476 75410
rect 164424 75346 164476 75352
rect 164436 21418 164464 75346
rect 164528 23118 164556 75886
rect 164620 75342 164648 79580
rect 164700 79562 164752 79568
rect 164700 79484 164752 79490
rect 164700 79426 164752 79432
rect 164712 75410 164740 79426
rect 164804 78946 164832 79784
rect 165034 79744 165062 80036
rect 164988 79716 165062 79744
rect 165126 79744 165154 80036
rect 165218 79812 165246 80036
rect 165310 79971 165338 80036
rect 165296 79962 165352 79971
rect 165296 79897 165352 79906
rect 165218 79784 165292 79812
rect 165126 79716 165200 79744
rect 164884 79620 164936 79626
rect 164884 79562 164936 79568
rect 164792 78940 164844 78946
rect 164792 78882 164844 78888
rect 164790 78704 164846 78713
rect 164790 78639 164846 78648
rect 164804 78402 164832 78639
rect 164792 78396 164844 78402
rect 164792 78338 164844 78344
rect 164792 77920 164844 77926
rect 164792 77862 164844 77868
rect 164700 75404 164752 75410
rect 164700 75346 164752 75352
rect 164608 75336 164660 75342
rect 164608 75278 164660 75284
rect 164700 75268 164752 75274
rect 164700 75210 164752 75216
rect 164608 75200 164660 75206
rect 164608 75142 164660 75148
rect 164516 23112 164568 23118
rect 164516 23054 164568 23060
rect 164620 23050 164648 75142
rect 164712 26926 164740 75210
rect 164804 57254 164832 77862
rect 164896 69834 164924 79562
rect 164988 75274 165016 79716
rect 165068 79484 165120 79490
rect 165068 79426 165120 79432
rect 165080 79286 165108 79426
rect 165068 79280 165120 79286
rect 165068 79222 165120 79228
rect 165068 79076 165120 79082
rect 165068 79018 165120 79024
rect 165080 78810 165108 79018
rect 165068 78804 165120 78810
rect 165068 78746 165120 78752
rect 165172 77926 165200 79716
rect 165160 77920 165212 77926
rect 165160 77862 165212 77868
rect 165066 77616 165122 77625
rect 165066 77551 165122 77560
rect 164976 75268 165028 75274
rect 164976 75210 165028 75216
rect 165080 72418 165108 77551
rect 165264 75914 165292 79784
rect 165402 79744 165430 80036
rect 165494 79812 165522 80036
rect 165586 79971 165614 80036
rect 165572 79962 165628 79971
rect 165572 79897 165628 79906
rect 165494 79784 165568 79812
rect 165402 79716 165476 79744
rect 165342 79656 165398 79665
rect 165342 79591 165398 79600
rect 165356 78198 165384 79591
rect 165448 78849 165476 79716
rect 165434 78840 165490 78849
rect 165434 78775 165490 78784
rect 165540 78577 165568 79784
rect 165678 79744 165706 80036
rect 165770 79966 165798 80036
rect 165862 79966 165890 80036
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165850 79960 165902 79966
rect 165850 79902 165902 79908
rect 165954 79898 165982 80036
rect 166046 79966 166074 80036
rect 166034 79960 166086 79966
rect 166034 79902 166086 79908
rect 165942 79892 165994 79898
rect 165942 79834 165994 79840
rect 166138 79830 166166 80036
rect 166034 79824 166086 79830
rect 166000 79772 166034 79778
rect 166000 79766 166086 79772
rect 166126 79824 166178 79830
rect 166230 79801 166258 80036
rect 166322 79966 166350 80036
rect 166310 79960 166362 79966
rect 166310 79902 166362 79908
rect 166414 79801 166442 80036
rect 166126 79766 166178 79772
rect 166216 79792 166272 79801
rect 165632 79716 165706 79744
rect 165804 79756 165856 79762
rect 165632 79014 165660 79716
rect 165804 79698 165856 79704
rect 166000 79750 166074 79766
rect 165710 79656 165766 79665
rect 165710 79591 165712 79600
rect 165764 79591 165766 79600
rect 165712 79562 165764 79568
rect 165620 79008 165672 79014
rect 165620 78950 165672 78956
rect 165712 78940 165764 78946
rect 165712 78882 165764 78888
rect 165618 78704 165674 78713
rect 165618 78639 165674 78648
rect 165526 78568 165582 78577
rect 165526 78503 165582 78512
rect 165344 78192 165396 78198
rect 165344 78134 165396 78140
rect 165172 75886 165292 75914
rect 165172 75206 165200 75886
rect 165160 75200 165212 75206
rect 165160 75142 165212 75148
rect 165068 72412 165120 72418
rect 165068 72354 165120 72360
rect 164884 69828 164936 69834
rect 164884 69770 164936 69776
rect 164792 57248 164844 57254
rect 164792 57190 164844 57196
rect 164700 26920 164752 26926
rect 164700 26862 164752 26868
rect 164608 23044 164660 23050
rect 164608 22986 164660 22992
rect 164424 21412 164476 21418
rect 164424 21354 164476 21360
rect 164332 14476 164384 14482
rect 164332 14418 164384 14424
rect 164240 7608 164292 7614
rect 164240 7550 164292 7556
rect 165632 4894 165660 78639
rect 165620 4888 165672 4894
rect 165620 4830 165672 4836
rect 165724 4826 165752 78882
rect 165816 78810 165844 79698
rect 165896 79688 165948 79694
rect 165896 79630 165948 79636
rect 165804 78804 165856 78810
rect 165804 78746 165856 78752
rect 165802 78704 165858 78713
rect 165802 78639 165858 78648
rect 165816 75410 165844 78639
rect 165804 75404 165856 75410
rect 165804 75346 165856 75352
rect 165804 75268 165856 75274
rect 165804 75210 165856 75216
rect 165816 11762 165844 75210
rect 165908 22982 165936 79630
rect 165896 22976 165948 22982
rect 165896 22918 165948 22924
rect 166000 22914 166028 79750
rect 166216 79727 166272 79736
rect 166400 79792 166456 79801
rect 166400 79727 166456 79736
rect 166172 79688 166224 79694
rect 166356 79688 166408 79694
rect 166172 79630 166224 79636
rect 166262 79656 166318 79665
rect 166080 79620 166132 79626
rect 166080 79562 166132 79568
rect 166092 78946 166120 79562
rect 166080 78940 166132 78946
rect 166080 78882 166132 78888
rect 166080 78804 166132 78810
rect 166080 78746 166132 78752
rect 166092 25770 166120 78746
rect 166184 29714 166212 79630
rect 166506 79676 166534 80036
rect 166598 79744 166626 80036
rect 166690 79937 166718 80036
rect 166676 79928 166732 79937
rect 166676 79863 166732 79872
rect 166782 79812 166810 80036
rect 166736 79784 166810 79812
rect 166598 79716 166672 79744
rect 166356 79630 166408 79636
rect 166460 79648 166534 79676
rect 166262 79591 166318 79600
rect 166276 31074 166304 79591
rect 166368 75274 166396 79630
rect 166356 75268 166408 75274
rect 166356 75210 166408 75216
rect 166460 70394 166488 79648
rect 166644 79626 166672 79716
rect 166632 79620 166684 79626
rect 166632 79562 166684 79568
rect 166540 79552 166592 79558
rect 166540 79494 166592 79500
rect 166552 79150 166580 79494
rect 166632 79348 166684 79354
rect 166632 79290 166684 79296
rect 166540 79144 166592 79150
rect 166540 79086 166592 79092
rect 166540 79008 166592 79014
rect 166540 78950 166592 78956
rect 166552 78742 166580 78950
rect 166644 78878 166672 79290
rect 166632 78872 166684 78878
rect 166632 78814 166684 78820
rect 166540 78736 166592 78742
rect 166736 78713 166764 79784
rect 166874 79744 166902 80036
rect 166966 79898 166994 80036
rect 166954 79892 167006 79898
rect 166954 79834 167006 79840
rect 167058 79778 167086 80036
rect 167150 79898 167178 80036
rect 167138 79892 167190 79898
rect 167138 79834 167190 79840
rect 166828 79716 166902 79744
rect 167012 79750 167086 79778
rect 167242 79778 167270 80036
rect 167334 79937 167362 80036
rect 167426 79966 167454 80036
rect 167414 79960 167466 79966
rect 167320 79928 167376 79937
rect 167414 79902 167466 79908
rect 167320 79863 167376 79872
rect 167368 79824 167420 79830
rect 167242 79750 167316 79778
rect 167518 79812 167546 80036
rect 167368 79766 167420 79772
rect 167472 79784 167546 79812
rect 166540 78678 166592 78684
rect 166722 78704 166778 78713
rect 166722 78639 166778 78648
rect 166630 78160 166686 78169
rect 166630 78095 166686 78104
rect 166644 77761 166672 78095
rect 166630 77752 166686 77761
rect 166630 77687 166686 77696
rect 166828 77625 166856 79716
rect 166906 79656 166962 79665
rect 166906 79591 166908 79600
rect 166960 79591 166962 79600
rect 166908 79562 166960 79568
rect 167012 79540 167040 79750
rect 167184 79688 167236 79694
rect 167184 79630 167236 79636
rect 167012 79512 167132 79540
rect 167000 79348 167052 79354
rect 167000 79290 167052 79296
rect 166908 79144 166960 79150
rect 166908 79086 166960 79092
rect 166920 78538 166948 79086
rect 167012 79014 167040 79290
rect 167000 79008 167052 79014
rect 167000 78950 167052 78956
rect 167000 78872 167052 78878
rect 167000 78814 167052 78820
rect 166908 78532 166960 78538
rect 166908 78474 166960 78480
rect 167012 78402 167040 78814
rect 167104 78402 167132 79512
rect 167000 78396 167052 78402
rect 167000 78338 167052 78344
rect 167092 78396 167144 78402
rect 167092 78338 167144 78344
rect 167090 78160 167146 78169
rect 167012 78118 167090 78146
rect 166814 77616 166870 77625
rect 166814 77551 166870 77560
rect 166724 75608 166776 75614
rect 166724 75550 166776 75556
rect 166736 75460 166764 75550
rect 166816 75472 166868 75478
rect 166736 75432 166816 75460
rect 166816 75414 166868 75420
rect 166540 75404 166592 75410
rect 166540 75346 166592 75352
rect 166368 70366 166488 70394
rect 166368 61402 166396 70366
rect 166552 69766 166580 75346
rect 167012 74526 167040 78118
rect 167090 78095 167146 78104
rect 167092 75132 167144 75138
rect 167092 75074 167144 75080
rect 167000 74520 167052 74526
rect 167000 74462 167052 74468
rect 166540 69760 166592 69766
rect 166540 69702 166592 69708
rect 166356 61396 166408 61402
rect 166356 61338 166408 61344
rect 166264 31068 166316 31074
rect 166264 31010 166316 31016
rect 166172 29708 166224 29714
rect 166172 29650 166224 29656
rect 166080 25764 166132 25770
rect 166080 25706 166132 25712
rect 165988 22908 166040 22914
rect 165988 22850 166040 22856
rect 167104 17270 167132 75074
rect 167196 24206 167224 79630
rect 167288 24274 167316 79750
rect 167380 24342 167408 79766
rect 167472 79676 167500 79784
rect 167610 79744 167638 80036
rect 167702 79937 167730 80036
rect 167688 79928 167744 79937
rect 167688 79863 167744 79872
rect 167794 79744 167822 80036
rect 167886 79937 167914 80036
rect 167872 79928 167928 79937
rect 167872 79863 167928 79872
rect 167610 79716 167684 79744
rect 167794 79716 167868 79744
rect 167472 79648 167592 79676
rect 167460 79348 167512 79354
rect 167460 79290 167512 79296
rect 167472 77518 167500 79290
rect 167460 77512 167512 77518
rect 167460 77454 167512 77460
rect 167460 75200 167512 75206
rect 167460 75142 167512 75148
rect 167472 29646 167500 75142
rect 167564 32502 167592 79648
rect 167656 78656 167684 79716
rect 167656 78628 167776 78656
rect 167642 78568 167698 78577
rect 167642 78503 167698 78512
rect 167656 66910 167684 78503
rect 167748 66978 167776 78628
rect 167840 75206 167868 79716
rect 167978 79676 168006 80036
rect 168070 79966 168098 80036
rect 168058 79960 168110 79966
rect 168058 79902 168110 79908
rect 168162 79898 168190 80036
rect 168254 79937 168282 80036
rect 168346 79966 168374 80036
rect 168334 79960 168386 79966
rect 168240 79928 168296 79937
rect 168150 79892 168202 79898
rect 168438 79937 168466 80036
rect 168334 79902 168386 79908
rect 168424 79928 168480 79937
rect 168240 79863 168296 79872
rect 168530 79898 168558 80036
rect 168622 79898 168650 80036
rect 168714 79898 168742 80036
rect 168806 79971 168834 80036
rect 168792 79962 168848 79971
rect 168424 79863 168480 79872
rect 168518 79892 168570 79898
rect 168150 79834 168202 79840
rect 168518 79834 168570 79840
rect 168610 79892 168662 79898
rect 168610 79834 168662 79840
rect 168702 79892 168754 79898
rect 168792 79897 168848 79906
rect 168702 79834 168754 79840
rect 168898 79812 168926 80036
rect 168990 79937 169018 80036
rect 168976 79928 169032 79937
rect 168976 79863 169032 79872
rect 169082 79812 169110 80036
rect 168852 79801 168926 79812
rect 169036 79801 169110 79812
rect 168562 79792 168618 79801
rect 168380 79756 168432 79762
rect 168380 79698 168432 79704
rect 168472 79756 168524 79762
rect 168562 79727 168618 79736
rect 168838 79792 168926 79801
rect 168894 79784 168926 79792
rect 169022 79792 169110 79801
rect 168838 79727 168894 79736
rect 169078 79784 169110 79792
rect 169174 79744 169202 80036
rect 169022 79727 169078 79736
rect 168472 79698 168524 79704
rect 168104 79688 168156 79694
rect 167978 79648 168052 79676
rect 168024 78792 168052 79648
rect 168104 79630 168156 79636
rect 168196 79688 168248 79694
rect 168196 79630 168248 79636
rect 167932 78764 168052 78792
rect 167828 75200 167880 75206
rect 167828 75142 167880 75148
rect 167932 75138 167960 78764
rect 168010 78704 168066 78713
rect 168010 78639 168066 78648
rect 167920 75132 167972 75138
rect 167920 75074 167972 75080
rect 168024 70394 168052 78639
rect 168116 77625 168144 79630
rect 168208 78169 168236 79630
rect 168288 78804 168340 78810
rect 168288 78746 168340 78752
rect 168194 78160 168250 78169
rect 168194 78095 168250 78104
rect 168102 77616 168158 77625
rect 168102 77551 168158 77560
rect 168300 77518 168328 78746
rect 168288 77512 168340 77518
rect 168288 77454 168340 77460
rect 168392 75206 168420 79698
rect 168380 75200 168432 75206
rect 168380 75142 168432 75148
rect 168380 75064 168432 75070
rect 168380 75006 168432 75012
rect 167932 70366 168052 70394
rect 167736 66972 167788 66978
rect 167736 66914 167788 66920
rect 167644 66904 167696 66910
rect 167644 66846 167696 66852
rect 167552 32496 167604 32502
rect 167552 32438 167604 32444
rect 167460 29640 167512 29646
rect 167460 29582 167512 29588
rect 167368 24336 167420 24342
rect 167368 24278 167420 24284
rect 167276 24268 167328 24274
rect 167276 24210 167328 24216
rect 167184 24200 167236 24206
rect 167184 24142 167236 24148
rect 167092 17264 167144 17270
rect 167092 17206 167144 17212
rect 167932 15910 167960 70366
rect 168392 18698 168420 75006
rect 168484 18766 168512 79698
rect 168576 75070 168604 79727
rect 169128 79716 169202 79744
rect 168656 79688 168708 79694
rect 168656 79630 168708 79636
rect 169024 79688 169076 79694
rect 169024 79630 169076 79636
rect 168668 78742 168696 79630
rect 168748 79552 168800 79558
rect 168748 79494 168800 79500
rect 168656 78736 168708 78742
rect 168656 78678 168708 78684
rect 168760 78441 168788 79494
rect 169036 78928 169064 79630
rect 168944 78900 169064 78928
rect 168944 78792 168972 78900
rect 168852 78764 168972 78792
rect 168746 78432 168802 78441
rect 168746 78367 168802 78376
rect 168748 78192 168800 78198
rect 168654 78160 168710 78169
rect 168748 78134 168800 78140
rect 168654 78095 168710 78104
rect 168564 75064 168616 75070
rect 168564 75006 168616 75012
rect 168564 74928 168616 74934
rect 168564 74870 168616 74876
rect 168472 18760 168524 18766
rect 168472 18702 168524 18708
rect 168380 18692 168432 18698
rect 168380 18634 168432 18640
rect 168576 18630 168604 74870
rect 168668 22846 168696 78095
rect 168760 77994 168788 78134
rect 168748 77988 168800 77994
rect 168748 77930 168800 77936
rect 168852 76537 168880 78764
rect 168930 78160 168986 78169
rect 168930 78095 168986 78104
rect 168838 76528 168894 76537
rect 168838 76463 168894 76472
rect 168748 75200 168800 75206
rect 168748 75142 168800 75148
rect 168840 75200 168892 75206
rect 168840 75142 168892 75148
rect 168760 24138 168788 75142
rect 168852 25634 168880 75142
rect 168944 62830 168972 78095
rect 169128 74934 169156 79716
rect 169266 79608 169294 80036
rect 169358 79676 169386 80036
rect 169450 79937 169478 80036
rect 169542 79966 169570 80036
rect 169530 79960 169582 79966
rect 169436 79928 169492 79937
rect 169634 79937 169662 80036
rect 169530 79902 169582 79908
rect 169620 79928 169676 79937
rect 169436 79863 169492 79872
rect 169620 79863 169676 79872
rect 169726 79812 169754 80036
rect 169680 79784 169754 79812
rect 169484 79688 169536 79694
rect 169358 79648 169432 79676
rect 169220 79580 169294 79608
rect 169116 74928 169168 74934
rect 169116 74870 169168 74876
rect 169220 70394 169248 79580
rect 169404 75206 169432 79648
rect 169484 79630 169536 79636
rect 169392 75200 169444 75206
rect 169392 75142 169444 75148
rect 169036 70366 169248 70394
rect 169036 64190 169064 70366
rect 169496 68338 169524 79630
rect 169574 78568 169630 78577
rect 169574 78503 169630 78512
rect 169588 75002 169616 78503
rect 169680 78169 169708 79784
rect 169818 79744 169846 80036
rect 169910 79971 169938 80036
rect 169896 79962 169952 79971
rect 169896 79897 169952 79906
rect 170002 79898 170030 80036
rect 170094 79971 170122 80036
rect 170080 79962 170136 79971
rect 169990 79892 170042 79898
rect 170080 79897 170136 79906
rect 169990 79834 170042 79840
rect 170186 79778 170214 80036
rect 170278 79937 170306 80036
rect 170264 79928 170320 79937
rect 170370 79898 170398 80036
rect 170462 79937 170490 80036
rect 170448 79928 170504 79937
rect 170264 79863 170320 79872
rect 170358 79892 170410 79898
rect 170448 79863 170504 79872
rect 170358 79834 170410 79840
rect 170554 79812 170582 80036
rect 170140 79750 170214 79778
rect 170508 79784 170582 79812
rect 170140 79744 170168 79750
rect 169772 79716 169846 79744
rect 170048 79716 170168 79744
rect 169666 78160 169722 78169
rect 169666 78095 169722 78104
rect 169772 75206 169800 79716
rect 169944 79688 169996 79694
rect 169944 79630 169996 79636
rect 169850 78704 169906 78713
rect 169850 78639 169906 78648
rect 169760 75200 169812 75206
rect 169760 75142 169812 75148
rect 169760 75064 169812 75070
rect 169760 75006 169812 75012
rect 169576 74996 169628 75002
rect 169576 74938 169628 74944
rect 169484 68332 169536 68338
rect 169484 68274 169536 68280
rect 169024 64184 169076 64190
rect 169024 64126 169076 64132
rect 168932 62824 168984 62830
rect 168932 62766 168984 62772
rect 168840 25628 168892 25634
rect 168840 25570 168892 25576
rect 168748 24132 168800 24138
rect 168748 24074 168800 24080
rect 168656 22840 168708 22846
rect 168656 22782 168708 22788
rect 168564 18624 168616 18630
rect 168564 18566 168616 18572
rect 167920 15904 167972 15910
rect 167920 15846 167972 15852
rect 165804 11756 165856 11762
rect 165804 11698 165856 11704
rect 169772 6186 169800 75006
rect 169864 6254 169892 78639
rect 169956 8974 169984 79630
rect 170048 25566 170076 79716
rect 170508 79665 170536 79784
rect 170646 79694 170674 80036
rect 170738 79937 170766 80036
rect 170724 79928 170780 79937
rect 170830 79898 170858 80036
rect 170922 79937 170950 80036
rect 170908 79928 170964 79937
rect 170724 79863 170780 79872
rect 170818 79892 170870 79898
rect 170908 79863 170964 79872
rect 170818 79834 170870 79840
rect 170726 79824 170778 79830
rect 170726 79766 170778 79772
rect 170634 79688 170686 79694
rect 170126 79656 170182 79665
rect 170126 79591 170182 79600
rect 170310 79656 170366 79665
rect 170310 79591 170366 79600
rect 170494 79656 170550 79665
rect 170634 79630 170686 79636
rect 170494 79591 170550 79600
rect 170140 78198 170168 79591
rect 170128 78192 170180 78198
rect 170128 78134 170180 78140
rect 170218 78160 170274 78169
rect 170218 78095 170274 78104
rect 170232 77897 170260 78095
rect 170218 77888 170274 77897
rect 170218 77823 170274 77832
rect 170324 77294 170352 79591
rect 170738 79540 170766 79766
rect 170864 79756 170916 79762
rect 171014 79744 171042 80036
rect 171106 79966 171134 80036
rect 171094 79960 171146 79966
rect 171198 79937 171226 80036
rect 171290 79966 171318 80036
rect 171278 79960 171330 79966
rect 171094 79902 171146 79908
rect 171184 79928 171240 79937
rect 171278 79902 171330 79908
rect 171184 79863 171240 79872
rect 171382 79830 171410 80036
rect 171474 79971 171502 80036
rect 171460 79962 171516 79971
rect 171460 79897 171516 79906
rect 171566 79898 171594 80036
rect 171658 79937 171686 80036
rect 171644 79928 171700 79937
rect 171554 79892 171606 79898
rect 171750 79898 171778 80036
rect 171644 79863 171700 79872
rect 171738 79892 171790 79898
rect 171554 79834 171606 79840
rect 171738 79834 171790 79840
rect 171232 79824 171284 79830
rect 171232 79766 171284 79772
rect 171370 79824 171422 79830
rect 171370 79766 171422 79772
rect 171598 79792 171654 79801
rect 170864 79698 170916 79704
rect 170968 79716 171042 79744
rect 170600 79512 170766 79540
rect 170496 78804 170548 78810
rect 170496 78746 170548 78752
rect 170324 77266 170444 77294
rect 170218 77072 170274 77081
rect 170218 77007 170274 77016
rect 170232 76673 170260 77007
rect 170218 76664 170274 76673
rect 170218 76599 170274 76608
rect 170416 75834 170444 77266
rect 170140 75806 170444 75834
rect 170140 32434 170168 75806
rect 170312 75200 170364 75206
rect 170312 75142 170364 75148
rect 170220 75132 170272 75138
rect 170220 75074 170272 75080
rect 170232 69018 170260 75074
rect 170324 69698 170352 75142
rect 170508 75070 170536 78746
rect 170600 78713 170628 79512
rect 170876 78810 170904 79698
rect 170864 78804 170916 78810
rect 170864 78746 170916 78752
rect 170586 78704 170642 78713
rect 170586 78639 170642 78648
rect 170862 78704 170918 78713
rect 170862 78639 170864 78648
rect 170916 78639 170918 78648
rect 170864 78610 170916 78616
rect 170862 78568 170918 78577
rect 170862 78503 170918 78512
rect 170680 78192 170732 78198
rect 170680 78134 170732 78140
rect 170496 75064 170548 75070
rect 170496 75006 170548 75012
rect 170312 69692 170364 69698
rect 170312 69634 170364 69640
rect 170220 69012 170272 69018
rect 170220 68954 170272 68960
rect 170128 32428 170180 32434
rect 170128 32370 170180 32376
rect 170692 25702 170720 78134
rect 170876 75138 170904 78503
rect 170864 75132 170916 75138
rect 170864 75074 170916 75080
rect 170968 73166 170996 79716
rect 171140 79688 171192 79694
rect 171046 79656 171102 79665
rect 171140 79630 171192 79636
rect 171046 79591 171102 79600
rect 171060 78198 171088 79591
rect 171048 78192 171100 78198
rect 171048 78134 171100 78140
rect 171152 75993 171180 79630
rect 171244 78470 171272 79766
rect 171508 79756 171560 79762
rect 171842 79744 171870 80036
rect 171598 79727 171654 79736
rect 171508 79698 171560 79704
rect 171520 79665 171548 79698
rect 171612 79694 171640 79727
rect 171704 79716 171870 79744
rect 171600 79688 171652 79694
rect 171506 79656 171562 79665
rect 171600 79630 171652 79636
rect 171506 79591 171562 79600
rect 171508 79552 171560 79558
rect 171508 79494 171560 79500
rect 171324 79008 171376 79014
rect 171324 78950 171376 78956
rect 171232 78464 171284 78470
rect 171232 78406 171284 78412
rect 171336 77450 171364 78950
rect 171520 78441 171548 79494
rect 171704 79098 171732 79716
rect 171934 79540 171962 80036
rect 172026 79642 172054 80036
rect 172118 79744 172146 80036
rect 172210 79812 172238 80036
rect 172302 79937 172330 80036
rect 172394 79966 172422 80036
rect 172382 79960 172434 79966
rect 172288 79928 172344 79937
rect 172486 79937 172514 80036
rect 172382 79902 172434 79908
rect 172472 79928 172528 79937
rect 172288 79863 172344 79872
rect 172578 79898 172606 80036
rect 172670 79898 172698 80036
rect 172472 79863 172528 79872
rect 172566 79892 172618 79898
rect 172566 79834 172618 79840
rect 172658 79892 172710 79898
rect 172658 79834 172710 79840
rect 172336 79824 172388 79830
rect 172210 79784 172284 79812
rect 172118 79716 172192 79744
rect 172026 79614 172100 79642
rect 171934 79512 172008 79540
rect 171784 79416 171836 79422
rect 171784 79358 171836 79364
rect 171612 79070 171732 79098
rect 171506 78432 171562 78441
rect 171506 78367 171562 78376
rect 171416 77648 171468 77654
rect 171416 77590 171468 77596
rect 171324 77444 171376 77450
rect 171324 77386 171376 77392
rect 171138 75984 171194 75993
rect 171138 75919 171194 75928
rect 170956 73160 171008 73166
rect 170956 73102 171008 73108
rect 171428 70394 171456 77590
rect 171612 77586 171640 79070
rect 171692 79008 171744 79014
rect 171692 78950 171744 78956
rect 171704 78538 171732 78950
rect 171796 78810 171824 79358
rect 171876 78872 171928 78878
rect 171876 78814 171928 78820
rect 171784 78804 171836 78810
rect 171784 78746 171836 78752
rect 171782 78704 171838 78713
rect 171782 78639 171784 78648
rect 171836 78639 171838 78648
rect 171784 78610 171836 78616
rect 171692 78532 171744 78538
rect 171692 78474 171744 78480
rect 171888 78418 171916 78814
rect 171980 78674 172008 79512
rect 171968 78668 172020 78674
rect 171968 78610 172020 78616
rect 172072 78538 172100 79614
rect 172164 79506 172192 79716
rect 172256 79626 172284 79784
rect 172762 79801 172790 80036
rect 172336 79766 172388 79772
rect 172748 79792 172804 79801
rect 172244 79620 172296 79626
rect 172244 79562 172296 79568
rect 172164 79478 172284 79506
rect 172152 79416 172204 79422
rect 172152 79358 172204 79364
rect 172164 78713 172192 79358
rect 172150 78704 172206 78713
rect 172150 78639 172206 78648
rect 172256 78577 172284 79478
rect 172348 78713 172376 79766
rect 172520 79756 172572 79762
rect 172748 79727 172804 79736
rect 172854 79744 172882 80036
rect 172946 79898 172974 80036
rect 172934 79892 172986 79898
rect 172934 79834 172986 79840
rect 173038 79744 173066 80036
rect 172854 79716 172928 79744
rect 172520 79698 172572 79704
rect 172428 79484 172480 79490
rect 172428 79426 172480 79432
rect 172334 78704 172390 78713
rect 172334 78639 172390 78648
rect 172440 78606 172468 79426
rect 172532 78878 172560 79698
rect 172612 79620 172664 79626
rect 172612 79562 172664 79568
rect 172520 78872 172572 78878
rect 172520 78814 172572 78820
rect 172428 78600 172480 78606
rect 172242 78568 172298 78577
rect 172060 78532 172112 78538
rect 172428 78542 172480 78548
rect 172242 78503 172298 78512
rect 172060 78474 172112 78480
rect 171888 78390 172192 78418
rect 171600 77580 171652 77586
rect 171600 77522 171652 77528
rect 171784 77512 171836 77518
rect 171784 77454 171836 77460
rect 171692 77444 171744 77450
rect 171692 77386 171744 77392
rect 171428 70366 171640 70394
rect 171612 43450 171640 70366
rect 171704 69902 171732 77386
rect 171692 69896 171744 69902
rect 171692 69838 171744 69844
rect 171692 69012 171744 69018
rect 171692 68954 171744 68960
rect 171600 43444 171652 43450
rect 171600 43386 171652 43392
rect 171704 33114 171732 68954
rect 171692 33108 171744 33114
rect 171692 33050 171744 33056
rect 170680 25696 170732 25702
rect 170680 25638 170732 25644
rect 170036 25560 170088 25566
rect 170036 25502 170088 25508
rect 169944 8968 169996 8974
rect 169944 8910 169996 8916
rect 169852 6248 169904 6254
rect 169852 6190 169904 6196
rect 169760 6180 169812 6186
rect 169760 6122 169812 6128
rect 169576 5228 169628 5234
rect 169576 5170 169628 5176
rect 164884 4820 164936 4826
rect 164884 4762 164936 4768
rect 165712 4820 165764 4826
rect 165712 4762 165764 4768
rect 163964 3732 164016 3738
rect 163964 3674 164016 3680
rect 162872 3454 163728 3482
rect 163700 480 163728 3454
rect 164896 480 164924 4762
rect 168380 3800 168432 3806
rect 168380 3742 168432 3748
rect 167184 3596 167236 3602
rect 167184 3538 167236 3544
rect 166080 3528 166132 3534
rect 166080 3470 166132 3476
rect 166092 480 166120 3470
rect 167196 480 167224 3538
rect 168392 480 168420 3742
rect 169588 480 169616 5170
rect 171796 3602 171824 77454
rect 172060 77376 172112 77382
rect 171966 77344 172022 77353
rect 172060 77318 172112 77324
rect 171966 77279 172022 77288
rect 171874 77208 171930 77217
rect 171874 77143 171876 77152
rect 171928 77143 171930 77152
rect 171876 77114 171928 77120
rect 171876 72412 171928 72418
rect 171876 72354 171928 72360
rect 171888 3670 171916 72354
rect 171980 17474 172008 77279
rect 171968 17468 172020 17474
rect 171968 17410 172020 17416
rect 171968 5024 172020 5030
rect 171968 4966 172020 4972
rect 171876 3664 171928 3670
rect 171876 3606 171928 3612
rect 171784 3596 171836 3602
rect 171784 3538 171836 3544
rect 170772 3460 170824 3466
rect 170772 3402 170824 3408
rect 170784 480 170812 3402
rect 171980 480 172008 4966
rect 172072 3874 172100 77318
rect 172164 3942 172192 78390
rect 172334 78296 172390 78305
rect 172334 78231 172390 78240
rect 172242 78160 172298 78169
rect 172242 78095 172298 78104
rect 172256 37942 172284 78095
rect 172348 39370 172376 78231
rect 172428 77716 172480 77722
rect 172428 77658 172480 77664
rect 172440 40730 172468 77658
rect 172624 77110 172652 79562
rect 172704 79484 172756 79490
rect 172704 79426 172756 79432
rect 172716 78441 172744 79426
rect 172702 78432 172758 78441
rect 172702 78367 172758 78376
rect 172612 77104 172664 77110
rect 172612 77046 172664 77052
rect 172900 76430 172928 79716
rect 172992 79716 173066 79744
rect 172992 79529 173020 79716
rect 173130 79642 173158 80036
rect 173222 79898 173250 80036
rect 173314 79937 173342 80036
rect 173300 79928 173356 79937
rect 173210 79892 173262 79898
rect 173300 79863 173356 79872
rect 173210 79834 173262 79840
rect 173256 79756 173308 79762
rect 173256 79698 173308 79704
rect 173084 79614 173158 79642
rect 172978 79520 173034 79529
rect 172978 79455 173034 79464
rect 173084 78985 173112 79614
rect 173268 79121 173296 79698
rect 173406 79676 173434 80036
rect 173498 79778 173526 80036
rect 173590 79966 173618 80036
rect 173682 79966 173710 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173670 79960 173722 79966
rect 173774 79937 173802 80036
rect 173670 79902 173722 79908
rect 173760 79928 173816 79937
rect 173760 79863 173816 79872
rect 173670 79824 173722 79830
rect 173668 79792 173670 79801
rect 173722 79792 173724 79801
rect 173498 79750 173572 79778
rect 173360 79648 173434 79676
rect 173360 79257 173388 79648
rect 173346 79248 173402 79257
rect 173346 79183 173402 79192
rect 173544 79121 173572 79750
rect 173866 79744 173894 80036
rect 173958 79966 173986 80036
rect 173946 79960 173998 79966
rect 173946 79902 173998 79908
rect 174050 79744 174078 80036
rect 174142 79898 174170 80036
rect 174130 79892 174182 79898
rect 174234 79880 174262 80036
rect 174340 80022 174492 80050
rect 174234 79852 174400 79880
rect 174130 79834 174182 79840
rect 174266 79792 174322 79801
rect 173668 79727 173724 79736
rect 173820 79716 173894 79744
rect 174004 79716 174078 79744
rect 174176 79756 174228 79762
rect 173624 79688 173676 79694
rect 173624 79630 173676 79636
rect 173254 79112 173310 79121
rect 173254 79047 173310 79056
rect 173530 79112 173586 79121
rect 173530 79047 173586 79056
rect 173070 78976 173126 78985
rect 173070 78911 173126 78920
rect 173636 78606 173664 79630
rect 173820 79626 173848 79716
rect 173808 79620 173860 79626
rect 173808 79562 173860 79568
rect 173624 78600 173676 78606
rect 173624 78542 173676 78548
rect 173164 78396 173216 78402
rect 173164 78338 173216 78344
rect 172888 76424 172940 76430
rect 172888 76366 172940 76372
rect 172518 60072 172574 60081
rect 172518 60007 172574 60016
rect 172428 40724 172480 40730
rect 172428 40666 172480 40672
rect 172336 39364 172388 39370
rect 172336 39306 172388 39312
rect 172244 37936 172296 37942
rect 172244 37878 172296 37884
rect 172532 16574 172560 60007
rect 172532 16546 172744 16574
rect 172152 3936 172204 3942
rect 172152 3878 172204 3884
rect 172060 3868 172112 3874
rect 172060 3810 172112 3816
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 3534 173204 78338
rect 174004 78305 174032 79716
rect 174266 79727 174322 79736
rect 174176 79698 174228 79704
rect 174188 79286 174216 79698
rect 174176 79280 174228 79286
rect 174176 79222 174228 79228
rect 174280 79218 174308 79727
rect 174268 79212 174320 79218
rect 174268 79154 174320 79160
rect 173990 78296 174046 78305
rect 173990 78231 174046 78240
rect 174372 78010 174400 79852
rect 174188 77982 174400 78010
rect 173254 76664 173310 76673
rect 173254 76599 173310 76608
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173268 3330 173296 76599
rect 173898 75712 173954 75721
rect 173898 75647 173954 75656
rect 173348 74520 173400 74526
rect 173348 74462 173400 74468
rect 173360 3466 173388 74462
rect 173348 3460 173400 3466
rect 173348 3402 173400 3408
rect 173256 3324 173308 3330
rect 173256 3266 173308 3272
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 75647
rect 173992 75200 174044 75206
rect 173992 75142 174044 75148
rect 174004 23322 174032 75142
rect 174188 64874 174216 77982
rect 174464 75914 174492 80022
rect 174544 80028 174596 80034
rect 174544 79970 174596 79976
rect 174556 79393 174584 79970
rect 174740 79490 174768 80650
rect 176016 80572 176068 80578
rect 176016 80514 176068 80520
rect 175280 80436 175332 80442
rect 175280 80378 175332 80384
rect 175188 80096 175240 80102
rect 175188 80038 175240 80044
rect 174728 79484 174780 79490
rect 174728 79426 174780 79432
rect 174542 79384 174598 79393
rect 174542 79319 174598 79328
rect 175200 78470 175228 80038
rect 175292 79422 175320 80378
rect 176028 80170 176056 80514
rect 176108 80504 176160 80510
rect 176108 80446 176160 80452
rect 176120 80170 176148 80446
rect 178328 80209 178356 80815
rect 178314 80200 178370 80209
rect 176016 80164 176068 80170
rect 176016 80106 176068 80112
rect 176108 80164 176160 80170
rect 178314 80135 178370 80144
rect 176108 80106 176160 80112
rect 178420 80034 178448 80951
rect 178500 80776 178552 80782
rect 178500 80718 178552 80724
rect 178408 80028 178460 80034
rect 178408 79970 178460 79976
rect 178512 79665 178540 80718
rect 178498 79656 178554 79665
rect 178498 79591 178554 79600
rect 175280 79416 175332 79422
rect 175280 79358 175332 79364
rect 178040 79416 178092 79422
rect 178040 79358 178092 79364
rect 175188 78464 175240 78470
rect 175188 78406 175240 78412
rect 174544 77852 174596 77858
rect 174544 77794 174596 77800
rect 174372 75886 174492 75914
rect 174372 75206 174400 75886
rect 174360 75200 174412 75206
rect 174360 75142 174412 75148
rect 174096 64846 174216 64874
rect 174096 45558 174124 64846
rect 174084 45552 174136 45558
rect 174084 45494 174136 45500
rect 173992 23316 174044 23322
rect 173992 23258 174044 23264
rect 174556 15978 174584 77794
rect 175924 77784 175976 77790
rect 175924 77726 175976 77732
rect 175278 69592 175334 69601
rect 175278 69527 175334 69536
rect 175292 16574 175320 69527
rect 175292 16546 175504 16574
rect 174544 15972 174596 15978
rect 174544 15914 174596 15920
rect 175476 480 175504 16546
rect 175936 6458 175964 77726
rect 176658 75576 176714 75585
rect 176658 75511 176714 75520
rect 176672 11694 176700 75511
rect 176752 27328 176804 27334
rect 176752 27270 176804 27276
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 27270
rect 178052 16574 178080 79358
rect 178972 78606 179000 82078
rect 179420 79348 179472 79354
rect 179420 79290 179472 79296
rect 179432 78674 179460 79290
rect 179420 78668 179472 78674
rect 179420 78610 179472 78616
rect 178960 78600 179012 78606
rect 178960 78542 179012 78548
rect 178774 77344 178830 77353
rect 178774 77279 178830 77288
rect 178788 77246 178816 77279
rect 178776 77240 178828 77246
rect 178776 77182 178828 77188
rect 178682 72720 178738 72729
rect 178682 72655 178738 72664
rect 178052 16546 178632 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 175924 6452 175976 6458
rect 175924 6394 175976 6400
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3806 178724 72655
rect 179616 71738 179644 135487
rect 180076 81297 180104 151778
rect 180156 146940 180208 146946
rect 180156 146882 180208 146888
rect 180168 131170 180196 146882
rect 180156 131164 180208 131170
rect 180156 131106 180208 131112
rect 180812 124137 180840 231066
rect 189724 205692 189776 205698
rect 189724 205634 189776 205640
rect 188344 165640 188396 165646
rect 188344 165582 188396 165588
rect 181260 162920 181312 162926
rect 181260 162862 181312 162868
rect 181168 142112 181220 142118
rect 181168 142054 181220 142060
rect 180984 141704 181036 141710
rect 180984 141646 181036 141652
rect 180890 137592 180946 137601
rect 180890 137527 180946 137536
rect 180798 124128 180854 124137
rect 180798 124063 180854 124072
rect 180156 111852 180208 111858
rect 180156 111794 180208 111800
rect 180062 81288 180118 81297
rect 180062 81223 180118 81232
rect 180168 80374 180196 111794
rect 180156 80368 180208 80374
rect 180156 80310 180208 80316
rect 180064 77920 180116 77926
rect 180064 77862 180116 77868
rect 179604 71732 179656 71738
rect 179604 71674 179656 71680
rect 179420 27260 179472 27266
rect 179420 27202 179472 27208
rect 179432 16574 179460 27202
rect 179432 16546 180012 16574
rect 178684 3800 178736 3806
rect 178684 3742 178736 3748
rect 179984 3482 180012 16546
rect 180076 5030 180104 77862
rect 180800 46232 180852 46238
rect 180800 46174 180852 46180
rect 180812 16574 180840 46174
rect 180904 33046 180932 137527
rect 180996 116657 181024 141646
rect 181076 140344 181128 140350
rect 181076 140286 181128 140292
rect 180982 116648 181038 116657
rect 180982 116583 181038 116592
rect 181088 112169 181116 140286
rect 181180 115161 181208 142054
rect 181272 133113 181300 162862
rect 182916 162172 182968 162178
rect 182916 162114 182968 162120
rect 182640 144492 182692 144498
rect 182640 144434 182692 144440
rect 182548 144424 182600 144430
rect 182548 144366 182600 144372
rect 182272 144356 182324 144362
rect 182272 144298 182324 144304
rect 182180 139460 182232 139466
rect 182180 139402 182232 139408
rect 182192 134609 182220 139402
rect 182178 134600 182234 134609
rect 182178 134535 182234 134544
rect 181258 133104 181314 133113
rect 181258 133039 181314 133048
rect 182180 131164 182232 131170
rect 182180 131106 182232 131112
rect 181166 115152 181222 115161
rect 181166 115087 181222 115096
rect 182192 113665 182220 131106
rect 182284 122641 182312 144298
rect 182456 141636 182508 141642
rect 182456 141578 182508 141584
rect 182364 140208 182416 140214
rect 182364 140150 182416 140156
rect 182270 122632 182326 122641
rect 182270 122567 182326 122576
rect 182376 118153 182404 140150
rect 182468 119649 182496 141578
rect 182560 127129 182588 144366
rect 182652 128625 182680 144434
rect 182732 140276 182784 140282
rect 182732 140218 182784 140224
rect 182638 128616 182694 128625
rect 182638 128551 182694 128560
rect 182546 127120 182602 127129
rect 182546 127055 182602 127064
rect 182744 121145 182772 140218
rect 182928 130121 182956 162114
rect 182914 130112 182970 130121
rect 182914 130047 182970 130056
rect 182824 125656 182876 125662
rect 182824 125598 182876 125604
rect 182730 121136 182786 121145
rect 182730 121071 182786 121080
rect 182454 119640 182510 119649
rect 182454 119575 182510 119584
rect 182362 118144 182418 118153
rect 182362 118079 182418 118088
rect 182178 113656 182234 113665
rect 182178 113591 182234 113600
rect 181074 112160 181130 112169
rect 181074 112095 181130 112104
rect 182836 86737 182864 125598
rect 183284 111784 183336 111790
rect 183284 111726 183336 111732
rect 183296 110673 183324 111726
rect 183282 110664 183338 110673
rect 183282 110599 183338 110608
rect 183468 110424 183520 110430
rect 183468 110366 183520 110372
rect 183480 109177 183508 110366
rect 183466 109168 183522 109177
rect 183466 109103 183522 109112
rect 183376 108996 183428 109002
rect 183376 108938 183428 108944
rect 183388 107681 183416 108938
rect 183374 107672 183430 107681
rect 183374 107607 183430 107616
rect 183468 106276 183520 106282
rect 183468 106218 183520 106224
rect 183480 106185 183508 106218
rect 183466 106176 183522 106185
rect 183466 106111 183522 106120
rect 183468 104848 183520 104854
rect 183468 104790 183520 104796
rect 183480 104689 183508 104790
rect 183466 104680 183522 104689
rect 183466 104615 183522 104624
rect 183468 103488 183520 103494
rect 183468 103430 183520 103436
rect 183480 103193 183508 103430
rect 183466 103184 183522 103193
rect 183466 103119 183522 103128
rect 183468 102128 183520 102134
rect 183468 102070 183520 102076
rect 183480 101697 183508 102070
rect 183466 101688 183522 101697
rect 183466 101623 183522 101632
rect 183468 100700 183520 100706
rect 183468 100642 183520 100648
rect 183480 100201 183508 100642
rect 183466 100192 183522 100201
rect 183466 100127 183522 100136
rect 183468 99340 183520 99346
rect 183468 99282 183520 99288
rect 183480 98705 183508 99282
rect 183466 98696 183522 98705
rect 183466 98631 183522 98640
rect 183468 97980 183520 97986
rect 183468 97922 183520 97928
rect 183480 97209 183508 97922
rect 183466 97200 183522 97209
rect 183466 97135 183522 97144
rect 183192 96620 183244 96626
rect 183192 96562 183244 96568
rect 183204 95713 183232 96562
rect 183190 95704 183246 95713
rect 183190 95639 183246 95648
rect 183284 95192 183336 95198
rect 183284 95134 183336 95140
rect 183296 94217 183324 95134
rect 183282 94208 183338 94217
rect 183282 94143 183338 94152
rect 183284 93832 183336 93838
rect 183284 93774 183336 93780
rect 183296 92721 183324 93774
rect 183282 92712 183338 92721
rect 183282 92647 183338 92656
rect 183468 92472 183520 92478
rect 183468 92414 183520 92420
rect 183480 91225 183508 92414
rect 183466 91216 183522 91225
rect 183466 91151 183522 91160
rect 183466 89720 183522 89729
rect 183466 89655 183468 89664
rect 183520 89655 183522 89664
rect 183468 89626 183520 89632
rect 188356 88262 188384 165582
rect 189736 89690 189764 205634
rect 207032 198014 207060 230588
rect 236012 230574 236578 230602
rect 207020 198008 207072 198014
rect 207020 197950 207072 197956
rect 236012 196722 236040 230574
rect 266556 228478 266584 230588
rect 266544 228472 266596 228478
rect 266544 228414 266596 228420
rect 267004 228472 267056 228478
rect 267004 228414 267056 228420
rect 236000 196716 236052 196722
rect 236000 196658 236052 196664
rect 267016 195906 267044 228414
rect 296732 199442 296760 230588
rect 296720 199436 296772 199442
rect 296720 199378 296772 199384
rect 327092 196654 327120 230588
rect 356532 228478 356560 230588
rect 356520 228472 356572 228478
rect 356520 228414 356572 228420
rect 377312 227044 377364 227050
rect 377312 226986 377364 226992
rect 377324 220114 377352 226986
rect 384396 226908 384448 226914
rect 384396 226850 384448 226856
rect 384408 224670 384436 226850
rect 381544 224664 381596 224670
rect 381544 224606 381596 224612
rect 384396 224664 384448 224670
rect 384396 224606 384448 224612
rect 368940 220108 368992 220114
rect 368940 220050 368992 220056
rect 377312 220108 377364 220114
rect 377312 220050 377364 220056
rect 368952 214606 368980 220050
rect 381556 216714 381584 224606
rect 386524 219434 386552 230588
rect 392676 229832 392728 229838
rect 392676 229774 392728 229780
rect 390928 229560 390980 229566
rect 390928 229502 390980 229508
rect 390940 226914 390968 229502
rect 390928 226908 390980 226914
rect 390928 226850 390980 226856
rect 386432 219406 386552 219434
rect 380164 216708 380216 216714
rect 380164 216650 380216 216656
rect 381544 216708 381596 216714
rect 381544 216650 381596 216656
rect 358728 214600 358780 214606
rect 358728 214542 358780 214548
rect 368940 214600 368992 214606
rect 368940 214542 368992 214548
rect 358740 211818 358768 214542
rect 344100 211812 344152 211818
rect 344100 211754 344152 211760
rect 358728 211812 358780 211818
rect 358728 211754 358780 211760
rect 344112 207058 344140 211754
rect 380176 208418 380204 216650
rect 376760 208412 376812 208418
rect 376760 208354 376812 208360
rect 380164 208412 380216 208418
rect 380164 208354 380216 208360
rect 341524 207052 341576 207058
rect 341524 206994 341576 207000
rect 344100 207052 344152 207058
rect 344100 206994 344152 207000
rect 341536 198762 341564 206994
rect 374000 202292 374052 202298
rect 374000 202234 374052 202240
rect 374012 199442 374040 202234
rect 376772 201346 376800 208354
rect 377680 204944 377732 204950
rect 377680 204886 377732 204892
rect 377692 202298 377720 204886
rect 377680 202292 377732 202298
rect 377680 202234 377732 202240
rect 375380 201340 375432 201346
rect 375380 201282 375432 201288
rect 376760 201340 376812 201346
rect 376760 201282 376812 201288
rect 351184 199436 351236 199442
rect 351184 199378 351236 199384
rect 374000 199436 374052 199442
rect 374000 199378 374052 199384
rect 338764 198756 338816 198762
rect 338764 198698 338816 198704
rect 341524 198756 341576 198762
rect 341524 198698 341576 198704
rect 327080 196648 327132 196654
rect 327080 196590 327132 196596
rect 267004 195900 267056 195906
rect 267004 195842 267056 195848
rect 338776 187746 338804 198698
rect 336004 187740 336056 187746
rect 336004 187682 336056 187688
rect 338764 187740 338816 187746
rect 338764 187682 338816 187688
rect 336016 178022 336044 187682
rect 330024 178016 330076 178022
rect 330024 177958 330076 177964
rect 336004 178016 336056 178022
rect 336004 177958 336056 177964
rect 330036 174146 330064 177958
rect 327724 174140 327776 174146
rect 327724 174082 327776 174088
rect 330024 174140 330076 174146
rect 330024 174082 330076 174088
rect 327736 161498 327764 174082
rect 351196 169794 351224 199378
rect 375392 196518 375420 201282
rect 367100 196512 367152 196518
rect 367100 196454 367152 196460
rect 375380 196512 375432 196518
rect 375380 196454 375432 196460
rect 367112 191842 367140 196454
rect 386432 195974 386460 219406
rect 392584 209840 392636 209846
rect 392584 209782 392636 209788
rect 389180 207052 389232 207058
rect 389180 206994 389232 207000
rect 389192 204950 389220 206994
rect 389180 204944 389232 204950
rect 389180 204886 389232 204892
rect 386420 195968 386472 195974
rect 386420 195910 386472 195916
rect 367020 191814 367140 191842
rect 367020 190534 367048 191814
rect 362224 190528 362276 190534
rect 362224 190470 362276 190476
rect 367008 190528 367060 190534
rect 367008 190470 367060 190476
rect 362236 172514 362264 190470
rect 392596 183530 392624 209782
rect 392688 207058 392716 229774
rect 392676 207052 392728 207058
rect 392676 206994 392728 207000
rect 390560 183524 390612 183530
rect 390560 183466 390612 183472
rect 392584 183524 392636 183530
rect 392584 183466 392636 183472
rect 390572 178106 390600 183466
rect 390480 178078 390600 178106
rect 390480 175234 390508 178078
rect 385684 175228 385736 175234
rect 385684 175170 385736 175176
rect 390468 175228 390520 175234
rect 390468 175170 390520 175176
rect 359832 172508 359884 172514
rect 359832 172450 359884 172456
rect 362224 172508 362276 172514
rect 362224 172450 362276 172456
rect 346308 169788 346360 169794
rect 346308 169730 346360 169736
rect 351184 169788 351236 169794
rect 351184 169730 351236 169736
rect 346320 166122 346348 169730
rect 340144 166116 340196 166122
rect 340144 166058 340196 166064
rect 346308 166116 346360 166122
rect 346308 166058 346360 166064
rect 324320 161492 324372 161498
rect 324320 161434 324372 161440
rect 327724 161492 327776 161498
rect 327724 161434 327776 161440
rect 324332 158778 324360 161434
rect 319904 158772 319956 158778
rect 319904 158714 319956 158720
rect 324320 158772 324372 158778
rect 324320 158714 324372 158720
rect 319916 155242 319944 158714
rect 340156 155242 340184 166058
rect 359844 165374 359872 172450
rect 356704 165368 356756 165374
rect 356704 165310 356756 165316
rect 359832 165368 359884 165374
rect 359832 165310 359884 165316
rect 356716 155990 356744 165310
rect 385696 160138 385724 175170
rect 382280 160132 382332 160138
rect 382280 160074 382332 160080
rect 385684 160132 385736 160138
rect 385684 160074 385736 160080
rect 382292 157434 382320 160074
rect 382200 157406 382320 157434
rect 382200 155990 382228 157406
rect 356704 155984 356756 155990
rect 356704 155926 356756 155932
rect 382188 155984 382240 155990
rect 382188 155926 382240 155932
rect 353944 155916 353996 155922
rect 353944 155858 353996 155864
rect 374644 155916 374696 155922
rect 374644 155858 374696 155864
rect 303988 155236 304040 155242
rect 303988 155178 304040 155184
rect 319904 155236 319956 155242
rect 319904 155178 319956 155184
rect 322204 155236 322256 155242
rect 322204 155178 322256 155184
rect 340144 155236 340196 155242
rect 340144 155178 340196 155184
rect 304000 152862 304028 155178
rect 301504 152856 301556 152862
rect 301504 152798 301556 152804
rect 303988 152856 304040 152862
rect 303988 152798 304040 152804
rect 301516 140146 301544 152798
rect 301504 140140 301556 140146
rect 301504 140082 301556 140088
rect 322216 134570 322244 155178
rect 353956 144838 353984 155858
rect 374656 150482 374684 155858
rect 372620 150476 372672 150482
rect 372620 150418 372672 150424
rect 374644 150476 374696 150482
rect 374644 150418 374696 150424
rect 372632 146334 372660 150418
rect 371884 146328 371936 146334
rect 371884 146270 371936 146276
rect 372620 146328 372672 146334
rect 372620 146270 372672 146276
rect 350540 144832 350592 144838
rect 350540 144774 350592 144780
rect 353944 144832 353996 144838
rect 353944 144774 353996 144780
rect 350552 136678 350580 144774
rect 371896 139466 371924 146270
rect 369768 139460 369820 139466
rect 369768 139402 369820 139408
rect 371884 139460 371936 139466
rect 371884 139402 371936 139408
rect 369780 138038 369808 139402
rect 367744 138032 367796 138038
rect 367744 137974 367796 137980
rect 369768 138032 369820 138038
rect 369768 137974 369820 137980
rect 350540 136672 350592 136678
rect 350540 136614 350592 136620
rect 345664 136604 345716 136610
rect 345664 136546 345716 136552
rect 295984 134564 296036 134570
rect 295984 134506 296036 134512
rect 322204 134564 322256 134570
rect 322204 134506 322256 134512
rect 295996 117026 296024 134506
rect 345676 124234 345704 136546
rect 367756 131170 367784 137974
rect 365720 131164 365772 131170
rect 365720 131106 365772 131112
rect 367744 131164 367796 131170
rect 367744 131106 367796 131112
rect 365732 127770 365760 131106
rect 363604 127764 363656 127770
rect 363604 127706 363656 127712
rect 365720 127764 365772 127770
rect 365720 127706 365772 127712
rect 345664 124228 345716 124234
rect 345664 124170 345716 124176
rect 342260 124160 342312 124166
rect 342260 124102 342312 124108
rect 293224 117020 293276 117026
rect 293224 116962 293276 116968
rect 295984 117020 296036 117026
rect 295984 116962 296036 116968
rect 189724 89684 189776 89690
rect 189724 89626 189776 89632
rect 183468 88256 183520 88262
rect 183466 88224 183468 88233
rect 188344 88256 188396 88262
rect 183520 88224 183522 88233
rect 188344 88198 188396 88204
rect 183466 88159 183522 88168
rect 182822 86728 182878 86737
rect 182822 86663 182878 86672
rect 183468 85604 183520 85610
rect 183468 85546 183520 85552
rect 183480 85241 183508 85546
rect 183466 85232 183522 85241
rect 183466 85167 183522 85176
rect 182822 83736 182878 83745
rect 182822 83671 182878 83680
rect 182180 80436 182232 80442
rect 182180 80378 182232 80384
rect 180892 33040 180944 33046
rect 180892 32982 180944 32988
rect 180812 16546 181024 16574
rect 180064 5024 180116 5030
rect 180064 4966 180116 4972
rect 179984 3454 180288 3482
rect 180260 480 180288 3454
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 80378
rect 182836 46918 182864 83671
rect 183466 82240 183522 82249
rect 183466 82175 183522 82184
rect 183480 81462 183508 82175
rect 183468 81456 183520 81462
rect 183468 81398 183520 81404
rect 200120 80300 200172 80306
rect 200120 80242 200172 80248
rect 195980 79144 196032 79150
rect 195980 79086 196032 79092
rect 194598 74080 194654 74089
rect 194598 74015 194654 74024
rect 184940 68672 184992 68678
rect 184940 68614 184992 68620
rect 182824 46912 182876 46918
rect 182824 46854 182876 46860
rect 183560 27192 183612 27198
rect 183560 27134 183612 27140
rect 183572 16574 183600 27134
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11694 184980 68614
rect 189080 67448 189132 67454
rect 189080 67390 189132 67396
rect 185032 61532 185084 61538
rect 185032 61474 185084 61480
rect 184940 11688 184992 11694
rect 184940 11630 184992 11636
rect 185044 6914 185072 61474
rect 187700 34128 187752 34134
rect 187700 34070 187752 34076
rect 186320 28484 186372 28490
rect 186320 28426 186372 28432
rect 186332 16574 186360 28426
rect 187712 16574 187740 34070
rect 189092 16574 189120 67390
rect 193218 65512 193274 65521
rect 193218 65447 193274 65456
rect 190460 28552 190512 28558
rect 190460 28494 190512 28500
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 11688 186188 11694
rect 186136 11630 186188 11636
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11630
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 28494
rect 191838 19000 191894 19009
rect 191838 18935 191894 18944
rect 191852 16574 191880 18935
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 65447
rect 193310 28520 193366 28529
rect 193310 28455 193366 28464
rect 193324 16574 193352 28455
rect 194612 16574 194640 74015
rect 195992 16574 196020 79086
rect 197360 76492 197412 76498
rect 197360 76434 197412 76440
rect 197372 16574 197400 76434
rect 198740 34060 198792 34066
rect 198740 34002 198792 34008
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 34002
rect 200132 16574 200160 80242
rect 231860 80232 231912 80238
rect 231860 80174 231912 80180
rect 213920 79008 213972 79014
rect 213920 78950 213972 78956
rect 211804 77036 211856 77042
rect 211804 76978 211856 76984
rect 209780 74248 209832 74254
rect 209780 74190 209832 74196
rect 202880 65952 202932 65958
rect 202880 65894 202932 65900
rect 201500 33992 201552 33998
rect 201500 33934 201552 33940
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11694 201540 33934
rect 201592 28416 201644 28422
rect 201592 28358 201644 28364
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 28358
rect 202892 16574 202920 65894
rect 207020 65884 207072 65890
rect 207020 65826 207072 65832
rect 205640 33924 205692 33930
rect 205640 33866 205692 33872
rect 204260 30116 204312 30122
rect 204260 30058 204312 30064
rect 204272 16574 204300 30058
rect 205652 16574 205680 33866
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 65826
rect 208400 30048 208452 30054
rect 208400 29990 208452 29996
rect 208412 16574 208440 29990
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 74190
rect 209872 70100 209924 70106
rect 209872 70042 209924 70048
rect 209884 16574 209912 70042
rect 209884 16546 211016 16574
rect 210988 480 211016 16546
rect 211816 3262 211844 76978
rect 213932 16574 213960 78950
rect 226340 76968 226392 76974
rect 226340 76910 226392 76916
rect 216680 74180 216732 74186
rect 216680 74122 216732 74128
rect 215300 24608 215352 24614
rect 215300 24550 215352 24556
rect 213932 16546 214512 16574
rect 213366 10704 213422 10713
rect 213366 10639 213422 10648
rect 212172 3324 212224 3330
rect 212172 3266 212224 3272
rect 211804 3256 211856 3262
rect 211804 3198 211856 3204
rect 212184 480 212212 3266
rect 213380 480 213408 10639
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 24550
rect 216692 16574 216720 74122
rect 223580 74112 223632 74118
rect 223580 74054 223632 74060
rect 218060 68604 218112 68610
rect 218060 68546 218112 68552
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 68546
rect 220820 65816 220872 65822
rect 220820 65758 220872 65764
rect 218152 24540 218204 24546
rect 218152 24482 218204 24488
rect 218164 16574 218192 24482
rect 220832 16574 220860 65758
rect 222200 26036 222252 26042
rect 222200 25978 222252 25984
rect 222212 16574 222240 25978
rect 218164 16546 219296 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 220452 5160 220504 5166
rect 220452 5102 220504 5108
rect 220464 480 220492 5102
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 74054
rect 225144 7948 225196 7954
rect 225144 7890 225196 7896
rect 225156 480 225184 7890
rect 226352 480 226380 76910
rect 230478 73944 230534 73953
rect 230478 73879 230534 73888
rect 227718 59936 227774 59945
rect 227718 59871 227774 59880
rect 226430 34096 226486 34105
rect 226430 34031 226486 34040
rect 226444 16574 226472 34031
rect 227732 16574 227760 59871
rect 229098 28384 229154 28393
rect 229098 28319 229154 28328
rect 229112 16574 229140 28319
rect 230492 16574 230520 73879
rect 226444 16546 227576 16574
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 80174
rect 252560 80164 252612 80170
rect 252560 80106 252612 80112
rect 249800 79076 249852 79082
rect 249800 79018 249852 79024
rect 247684 78328 247736 78334
rect 247684 78270 247736 78276
rect 247038 76936 247094 76945
rect 240140 76900 240192 76906
rect 247038 76871 247094 76880
rect 240140 76842 240192 76848
rect 234620 64524 234672 64530
rect 234620 64466 234672 64472
rect 233240 29980 233292 29986
rect 233240 29922 233292 29928
rect 233252 16574 233280 29922
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 64466
rect 238760 64456 238812 64462
rect 238760 64398 238812 64404
rect 234712 33856 234764 33862
rect 234712 33798 234764 33804
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 33798
rect 236000 29912 236052 29918
rect 236000 29854 236052 29860
rect 236012 16574 236040 29854
rect 238772 16574 238800 64398
rect 236012 16546 236592 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 12028 237708 12034
rect 237656 11970 237708 11976
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 11970
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 76842
rect 244278 73808 244334 73817
rect 244278 73743 244334 73752
rect 242900 31476 242952 31482
rect 242900 31418 242952 31424
rect 241704 14816 241756 14822
rect 241704 14758 241756 14764
rect 241716 480 241744 14758
rect 242912 4214 242940 31418
rect 244292 16574 244320 73743
rect 247052 16574 247080 76871
rect 247696 20194 247724 78270
rect 248418 20224 248474 20233
rect 247684 20188 247736 20194
rect 248418 20159 248474 20168
rect 247684 20130 247736 20136
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 242992 7880 243044 7886
rect 242992 7822 243044 7828
rect 242900 4208 242952 4214
rect 242900 4150 242952 4156
rect 243004 3482 243032 7822
rect 244096 4208 244148 4214
rect 244096 4150 244148 4156
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 4150
rect 245212 480 245240 16546
rect 246394 7712 246450 7721
rect 246394 7647 246450 7656
rect 246408 480 246436 7647
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 20159
rect 249812 16574 249840 79018
rect 251180 74044 251232 74050
rect 251180 73986 251232 73992
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 4214 251220 73986
rect 251272 65748 251324 65754
rect 251272 65690 251324 65696
rect 251180 4208 251232 4214
rect 251180 4150 251232 4156
rect 251284 3482 251312 65690
rect 252572 16574 252600 80106
rect 267740 78940 267792 78946
rect 267740 78882 267792 78888
rect 253204 78260 253256 78266
rect 253204 78202 253256 78208
rect 253216 20126 253244 78202
rect 260840 76832 260892 76838
rect 260840 76774 260892 76780
rect 256700 65680 256752 65686
rect 256700 65622 256752 65628
rect 253940 29844 253992 29850
rect 253940 29786 253992 29792
rect 253204 20120 253256 20126
rect 253204 20062 253256 20068
rect 253952 16574 253980 29786
rect 255320 20392 255372 20398
rect 255320 20334 255372 20340
rect 255332 16574 255360 20334
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 4208 252428 4214
rect 252376 4150 252428 4156
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 4150
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 65622
rect 259460 35624 259512 35630
rect 259460 35566 259512 35572
rect 258080 29776 258132 29782
rect 258080 29718 258132 29724
rect 258092 16574 258120 29718
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 480 259500 35566
rect 260852 16574 260880 76774
rect 266358 33960 266414 33969
rect 266358 33895 266414 33904
rect 262220 20324 262272 20330
rect 262220 20266 262272 20272
rect 262232 16574 262260 20266
rect 266372 16574 266400 33895
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 260656 9308 260708 9314
rect 260656 9250 260708 9256
rect 260668 480 260696 9250
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264150 9208 264206 9217
rect 264150 9143 264206 9152
rect 264164 480 264192 9143
rect 265346 7576 265402 7585
rect 265346 7511 265402 7520
rect 265360 480 265388 7511
rect 266556 480 266584 16546
rect 267752 480 267780 78882
rect 293236 78878 293264 116962
rect 342272 116006 342300 124102
rect 363616 117706 363644 127706
rect 360200 117700 360252 117706
rect 360200 117642 360252 117648
rect 363604 117700 363656 117706
rect 363604 117642 363656 117648
rect 342260 116000 342312 116006
rect 342260 115942 342312 115948
rect 338764 115932 338816 115938
rect 338764 115874 338816 115880
rect 338776 111926 338804 115874
rect 360212 115122 360240 117642
rect 358268 115116 358320 115122
rect 358268 115058 358320 115064
rect 360200 115116 360252 115122
rect 360200 115058 360252 115064
rect 358280 113830 358308 115058
rect 351920 113824 351972 113830
rect 351920 113766 351972 113772
rect 358268 113824 358320 113830
rect 358268 113766 358320 113772
rect 351932 111926 351960 113766
rect 336740 111920 336792 111926
rect 336740 111862 336792 111868
rect 338764 111920 338816 111926
rect 338764 111862 338816 111868
rect 349160 111920 349212 111926
rect 349160 111862 349212 111868
rect 351920 111920 351972 111926
rect 351920 111862 351972 111868
rect 336752 111790 336780 111862
rect 336740 111784 336792 111790
rect 336740 111726 336792 111732
rect 349172 110498 349200 111862
rect 349160 110492 349212 110498
rect 349160 110434 349212 110440
rect 393976 80782 394004 231814
rect 394712 229566 394740 232086
rect 394700 229560 394752 229566
rect 394700 229502 394752 229508
rect 396460 220794 396488 678234
rect 396540 647216 396592 647222
rect 396540 647158 396592 647164
rect 396552 243574 396580 647158
rect 396724 643136 396776 643142
rect 396724 643078 396776 643084
rect 396632 536444 396684 536450
rect 396632 536386 396684 536392
rect 396540 243568 396592 243574
rect 396540 243510 396592 243516
rect 396540 240100 396592 240106
rect 396540 240042 396592 240048
rect 396552 238882 396580 240042
rect 396540 238876 396592 238882
rect 396540 238818 396592 238824
rect 396540 238740 396592 238746
rect 396540 238682 396592 238688
rect 396552 232150 396580 238682
rect 396540 232144 396592 232150
rect 396540 232086 396592 232092
rect 396540 232008 396592 232014
rect 396540 231950 396592 231956
rect 396552 227050 396580 231950
rect 396644 229838 396672 536386
rect 396632 229832 396684 229838
rect 396632 229774 396684 229780
rect 396540 227044 396592 227050
rect 396540 226986 396592 226992
rect 394056 220788 394108 220794
rect 394056 220730 394108 220736
rect 396448 220788 396500 220794
rect 396448 220730 396500 220736
rect 394068 209846 394096 220730
rect 394056 209840 394108 209846
rect 394056 209782 394108 209788
rect 393964 80776 394016 80782
rect 393964 80718 394016 80724
rect 293224 78872 293276 78878
rect 293224 78814 293276 78820
rect 396736 78577 396764 643078
rect 396816 378208 396868 378214
rect 396816 378150 396868 378156
rect 396828 81161 396856 378150
rect 397000 324352 397052 324358
rect 397000 324294 397052 324300
rect 396908 243568 396960 243574
rect 396908 243510 396960 243516
rect 396920 232014 396948 243510
rect 396908 232008 396960 232014
rect 396908 231950 396960 231956
rect 396814 81152 396870 81161
rect 396814 81087 396870 81096
rect 397012 81025 397040 324294
rect 396998 81016 397054 81025
rect 396998 80951 397054 80960
rect 397472 78849 397500 703520
rect 410524 700460 410576 700466
rect 410524 700402 410576 700408
rect 409144 700392 409196 700398
rect 409144 700334 409196 700340
rect 407764 700324 407816 700330
rect 407764 700266 407816 700272
rect 406384 670744 406436 670750
rect 406384 670686 406436 670692
rect 405004 616888 405056 616894
rect 405004 616830 405056 616836
rect 403624 563100 403676 563106
rect 403624 563042 403676 563048
rect 400864 510672 400916 510678
rect 400864 510614 400916 510620
rect 399484 456816 399536 456822
rect 399484 456758 399536 456764
rect 398104 418192 398156 418198
rect 398104 418134 398156 418140
rect 398116 144226 398144 418134
rect 398196 364404 398248 364410
rect 398196 364346 398248 364352
rect 398208 144294 398236 364346
rect 398288 311908 398340 311914
rect 398288 311850 398340 311856
rect 398196 144288 398248 144294
rect 398196 144230 398248 144236
rect 398104 144220 398156 144226
rect 398104 144162 398156 144168
rect 398300 142934 398328 311850
rect 398380 258120 398432 258126
rect 398380 258062 398432 258068
rect 398392 143002 398420 258062
rect 398380 142996 398432 143002
rect 398380 142938 398432 142944
rect 398288 142928 398340 142934
rect 398288 142870 398340 142876
rect 399496 97986 399524 456758
rect 400876 99346 400904 510614
rect 403636 100706 403664 563042
rect 405016 102134 405044 616830
rect 406396 103494 406424 670686
rect 407776 104854 407804 700266
rect 409156 106282 409184 700334
rect 410536 109002 410564 700402
rect 412652 140078 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 418804 404388 418856 404394
rect 418804 404330 418856 404336
rect 417424 351960 417476 351966
rect 417424 351902 417476 351908
rect 414664 298172 414716 298178
rect 414664 298114 414716 298120
rect 413284 244316 413336 244322
rect 413284 244258 413336 244264
rect 412640 140072 412692 140078
rect 412640 140014 412692 140020
rect 410524 108996 410576 109002
rect 410524 108938 410576 108944
rect 409144 106276 409196 106282
rect 409144 106218 409196 106224
rect 407764 104848 407816 104854
rect 407764 104790 407816 104796
rect 406384 103488 406436 103494
rect 406384 103430 406436 103436
rect 405004 102128 405056 102134
rect 405004 102070 405056 102076
rect 403624 100700 403676 100706
rect 403624 100642 403676 100648
rect 400864 99340 400916 99346
rect 400864 99282 400916 99288
rect 399484 97980 399536 97986
rect 399484 97922 399536 97928
rect 413296 92478 413324 244258
rect 414676 93838 414704 298114
rect 417436 95198 417464 351902
rect 418816 96626 418844 404330
rect 418804 96620 418856 96626
rect 418804 96562 418856 96568
rect 417424 95192 417476 95198
rect 417424 95134 417476 95140
rect 414664 93832 414716 93838
rect 414664 93774 414716 93780
rect 413284 92472 413336 92478
rect 413284 92414 413336 92420
rect 430580 80096 430632 80102
rect 430580 80038 430632 80044
rect 397458 78840 397514 78849
rect 397458 78775 397514 78784
rect 396722 78568 396778 78577
rect 396722 78503 396778 78512
rect 322204 78192 322256 78198
rect 322204 78134 322256 78140
rect 282918 76800 282974 76809
rect 282918 76735 282974 76744
rect 288440 76764 288492 76770
rect 270500 67380 270552 67386
rect 270500 67322 270552 67328
rect 269120 33788 269172 33794
rect 269120 33730 269172 33736
rect 267832 31408 267884 31414
rect 267832 31350 267884 31356
rect 267844 16574 267872 31350
rect 269132 16574 269160 33730
rect 270512 16574 270540 67322
rect 274640 63164 274692 63170
rect 274640 63106 274692 63112
rect 271880 28348 271932 28354
rect 271880 28290 271932 28296
rect 271892 16574 271920 28290
rect 273260 20256 273312 20262
rect 273260 20198 273312 20204
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 20198
rect 274652 16574 274680 63106
rect 280158 44840 280214 44849
rect 280158 44775 280214 44784
rect 276020 35556 276072 35562
rect 276020 35498 276072 35504
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 4214 276060 35498
rect 276112 27124 276164 27130
rect 276112 27066 276164 27072
rect 276020 4208 276072 4214
rect 276020 4150 276072 4156
rect 276124 3482 276152 27066
rect 278780 25968 278832 25974
rect 278780 25910 278832 25916
rect 278792 16574 278820 25910
rect 280172 16574 280200 44775
rect 282932 16574 282960 76735
rect 288440 76706 288492 76712
rect 284298 72584 284354 72593
rect 284298 72519 284354 72528
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 278320 9240 278372 9246
rect 278320 9182 278372 9188
rect 276756 4208 276808 4214
rect 276756 4150 276808 4156
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 4150
rect 278332 480 278360 9182
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281538 10568 281594 10577
rect 281538 10503 281594 10512
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 10503
rect 283116 480 283144 16546
rect 284312 480 284340 72519
rect 284392 71052 284444 71058
rect 284392 70994 284444 71000
rect 284404 16574 284432 70994
rect 287060 35488 287112 35494
rect 287060 35430 287112 35436
rect 285680 28280 285732 28286
rect 285680 28222 285732 28228
rect 285692 16574 285720 28222
rect 287072 16574 287100 35430
rect 288452 16574 288480 76706
rect 296720 76696 296772 76702
rect 296720 76638 296772 76644
rect 291200 72684 291252 72690
rect 291200 72626 291252 72632
rect 289820 31340 289872 31346
rect 289820 31282 289872 31288
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 31282
rect 291212 16574 291240 72626
rect 292580 64388 292632 64394
rect 292580 64330 292632 64336
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 64330
rect 293960 35420 294012 35426
rect 293960 35362 294012 35368
rect 292672 24472 292724 24478
rect 292672 24414 292724 24420
rect 292684 16574 292712 24414
rect 293972 16574 294000 35362
rect 296732 16574 296760 76638
rect 318800 73976 318852 73982
rect 318800 73918 318852 73924
rect 311900 72616 311952 72622
rect 311900 72558 311952 72564
rect 298098 72448 298154 72457
rect 298098 72383 298154 72392
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 295616 10600 295668 10606
rect 295616 10542 295668 10548
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 10542
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 72383
rect 306380 67312 306432 67318
rect 306380 67254 306432 67260
rect 305000 35352 305052 35358
rect 305000 35294 305052 35300
rect 303620 23384 303672 23390
rect 303620 23326 303672 23332
rect 303632 16574 303660 23326
rect 305012 16574 305040 35294
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301502 13288 301558 13297
rect 301502 13223 301558 13232
rect 299662 10432 299718 10441
rect 299662 10367 299718 10376
rect 299676 480 299704 10367
rect 300766 9072 300822 9081
rect 300766 9007 300822 9016
rect 300780 480 300808 9007
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 13223
rect 303160 3868 303212 3874
rect 303160 3810 303212 3816
rect 303172 480 303200 3810
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 67254
rect 309140 63096 309192 63102
rect 309140 63038 309192 63044
rect 307760 35284 307812 35290
rect 307760 35226 307812 35232
rect 307772 3262 307800 35226
rect 307852 25900 307904 25906
rect 307852 25842 307904 25848
rect 307864 16574 307892 25842
rect 309152 16574 309180 63038
rect 310520 27056 310572 27062
rect 310520 26998 310572 27004
rect 310532 16574 310560 26998
rect 311912 16574 311940 72558
rect 316038 53136 316094 53145
rect 316038 53071 316094 53080
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307760 3256 307812 3262
rect 307760 3198 307812 3204
rect 307956 480 307984 16546
rect 309048 3256 309100 3262
rect 309048 3198 309100 3204
rect 309060 480 309088 3198
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313832 11960 313884 11966
rect 313832 11902 313884 11908
rect 313844 480 313872 11902
rect 315026 5128 315082 5137
rect 315026 5063 315082 5072
rect 315040 480 315068 5063
rect 316052 3262 316080 53071
rect 317418 29608 317474 29617
rect 317418 29543 317474 29552
rect 317432 16574 317460 29543
rect 318812 16574 318840 73918
rect 320180 68536 320232 68542
rect 320180 68478 320232 68484
rect 319442 21720 319498 21729
rect 319442 21655 319498 21664
rect 317432 16546 318104 16574
rect 318812 16546 319392 16574
rect 316222 16280 316278 16289
rect 316222 16215 316278 16224
rect 316040 3256 316092 3262
rect 316040 3198 316092 3204
rect 316236 480 316264 16215
rect 317328 3256 317380 3262
rect 317328 3198 317380 3204
rect 317340 480 317368 3198
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319364 3482 319392 16546
rect 319456 3874 319484 21655
rect 320192 16574 320220 68478
rect 322216 28286 322244 78134
rect 324412 76628 324464 76634
rect 324412 76570 324464 76576
rect 322204 28280 322256 28286
rect 322204 28222 322256 28228
rect 320192 16546 320496 16574
rect 319444 3868 319496 3874
rect 319444 3810 319496 3816
rect 319364 3454 319760 3482
rect 319732 480 319760 3454
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 323308 6792 323360 6798
rect 323308 6734 323360 6740
rect 322112 3392 322164 3398
rect 322112 3334 322164 3340
rect 322124 480 322152 3334
rect 323320 480 323348 6734
rect 324424 480 324452 76570
rect 396080 75608 396132 75614
rect 396080 75550 396132 75556
rect 354680 73908 354732 73914
rect 354680 73850 354732 73856
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 338120 64320 338172 64326
rect 338120 64262 338172 64268
rect 332600 31272 332652 31278
rect 332600 31214 332652 31220
rect 332612 16574 332640 31214
rect 338132 16574 338160 64262
rect 339500 26988 339552 26994
rect 339500 26930 339552 26936
rect 332612 16546 332732 16574
rect 338132 16546 338712 16574
rect 326804 6724 326856 6730
rect 326804 6666 326856 6672
rect 325608 4140 325660 4146
rect 325608 4082 325660 4088
rect 325620 480 325648 4082
rect 326816 480 326844 6666
rect 329196 6656 329248 6662
rect 329196 6598 329248 6604
rect 328000 4072 328052 4078
rect 328000 4014 328052 4020
rect 328012 480 328040 4014
rect 329208 480 329236 6598
rect 330392 6588 330444 6594
rect 330392 6530 330444 6536
rect 330404 480 330432 6530
rect 331588 4004 331640 4010
rect 331588 3946 331640 3952
rect 331600 480 331628 3946
rect 332704 480 332732 16546
rect 336278 6488 336334 6497
rect 336278 6423 336334 6432
rect 333886 6216 333942 6225
rect 333886 6151 333942 6160
rect 333900 480 333928 6151
rect 335082 3632 335138 3641
rect 335082 3567 335138 3576
rect 335096 480 335124 3567
rect 336292 480 336320 6423
rect 337474 6352 337530 6361
rect 337474 6287 337530 6296
rect 337488 480 337516 6287
rect 338684 480 338712 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 26930
rect 340892 3210 340920 72490
rect 353298 71224 353354 71233
rect 353298 71159 353354 71168
rect 347780 67244 347832 67250
rect 347780 67186 347832 67192
rect 340972 67176 341024 67182
rect 340972 67118 341024 67124
rect 340984 3398 341012 67118
rect 346400 25832 346452 25838
rect 346400 25774 346452 25780
rect 343640 21684 343692 21690
rect 343640 21626 343692 21632
rect 343652 16574 343680 21626
rect 346412 16574 346440 25774
rect 347792 16574 347820 67186
rect 351918 47560 351974 47569
rect 351918 47495 351974 47504
rect 350538 18864 350594 18873
rect 350538 18799 350594 18808
rect 350552 16574 350580 18799
rect 351932 16574 351960 47495
rect 353312 16574 353340 71159
rect 354692 16574 354720 73850
rect 375380 73840 375432 73846
rect 375380 73782 375432 73788
rect 357440 72480 357492 72486
rect 357440 72422 357492 72428
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 343364 9172 343416 9178
rect 343364 9114 343416 9120
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 343376 480 343404 9114
rect 344572 480 344600 16546
rect 345296 13456 345348 13462
rect 345296 13398 345348 13404
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 13398
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349160 13388 349212 13394
rect 349160 13330 349212 13336
rect 349172 3210 349200 13330
rect 349250 13152 349306 13161
rect 349250 13087 349306 13096
rect 349264 3398 349292 13087
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356336 3936 356388 3942
rect 356336 3878 356388 3884
rect 356348 480 356376 3878
rect 357452 3398 357480 72422
rect 362960 68468 363012 68474
rect 362960 68410 363012 68416
rect 358820 65612 358872 65618
rect 358820 65554 358872 65560
rect 357532 31204 357584 31210
rect 357532 31146 357584 31152
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 31146
rect 358832 16574 358860 65554
rect 360200 23248 360252 23254
rect 360200 23190 360252 23196
rect 360212 16574 360240 23190
rect 362972 16574 363000 68410
rect 368480 64252 368532 64258
rect 368480 64194 368532 64200
rect 367098 40624 367154 40633
rect 367098 40559 367154 40568
rect 367112 16574 367140 40559
rect 368492 16574 368520 64194
rect 374000 63028 374052 63034
rect 374000 62970 374052 62976
rect 372618 35184 372674 35193
rect 372618 35119 372674 35128
rect 372632 16574 372660 35119
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 362972 16546 363552 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 372632 16546 372936 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 362316 3324 362368 3330
rect 362316 3266 362368 3272
rect 362328 480 362356 3266
rect 363524 480 363552 16546
rect 365720 13320 365772 13326
rect 365720 13262 365772 13268
rect 364616 10532 364668 10538
rect 364616 10474 364668 10480
rect 364628 480 364656 10474
rect 365732 3398 365760 13262
rect 365812 5092 365864 5098
rect 365812 5034 365864 5040
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 5034
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 371238 16144 371294 16153
rect 371238 16079 371294 16088
rect 370134 14784 370190 14793
rect 370134 14719 370190 14728
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 14719
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 16079
rect 372908 480 372936 16546
rect 374012 1170 374040 62970
rect 374092 24404 374144 24410
rect 374092 24346 374144 24352
rect 374104 3398 374132 24346
rect 375392 16574 375420 73782
rect 382280 70032 382332 70038
rect 382280 69974 382332 69980
rect 376760 65544 376812 65550
rect 376760 65486 376812 65492
rect 376772 16574 376800 65486
rect 379520 23180 379572 23186
rect 379520 23122 379572 23128
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378416 16176 378468 16182
rect 378416 16118 378468 16124
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16118
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 23122
rect 381176 14748 381228 14754
rect 381176 14690 381228 14696
rect 381188 480 381216 14690
rect 382292 3210 382320 69974
rect 390560 69964 390612 69970
rect 390560 69906 390612 69912
rect 382372 35216 382424 35222
rect 382372 35158 382424 35164
rect 382384 3398 382412 35158
rect 389180 31136 389232 31142
rect 389180 31078 389232 31084
rect 386418 25528 386474 25537
rect 386418 25463 386474 25472
rect 386432 16574 386460 25463
rect 389192 16574 389220 31078
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 384304 14680 384356 14686
rect 384304 14622 384356 14628
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14622
rect 385960 14612 386012 14618
rect 385960 14554 386012 14560
rect 385972 480 386000 14554
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387798 16008 387854 16017
rect 387798 15943 387854 15952
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 15943
rect 389468 480 389496 16546
rect 390572 1290 390600 69906
rect 390652 42084 390704 42090
rect 390652 42026 390704 42032
rect 390560 1284 390612 1290
rect 390560 1226 390612 1232
rect 390664 480 390692 42026
rect 391940 32768 391992 32774
rect 391940 32710 391992 32716
rect 391952 16574 391980 32710
rect 391952 16546 392624 16574
rect 391848 1284 391900 1290
rect 391848 1226 391900 1232
rect 391860 480 391888 1226
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 395344 16108 395396 16114
rect 395344 16050 395396 16056
rect 394240 10464 394292 10470
rect 394240 10406 394292 10412
rect 394252 480 394280 10406
rect 395356 480 395384 16050
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 75550
rect 402978 75440 403034 75449
rect 402978 75375 403034 75384
rect 401600 58676 401652 58682
rect 401600 58618 401652 58624
rect 397460 37936 397512 37942
rect 397460 37878 397512 37884
rect 397472 16574 397500 37878
rect 401612 16574 401640 58618
rect 402992 16574 403020 75375
rect 426440 69896 426492 69902
rect 426440 69838 426492 69844
rect 408500 62960 408552 62966
rect 408500 62902 408552 62908
rect 404360 39364 404412 39370
rect 404360 39306 404412 39312
rect 397472 16546 397776 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 397748 480 397776 16546
rect 398840 16040 398892 16046
rect 398840 15982 398892 15988
rect 398852 3210 398880 15982
rect 398932 10396 398984 10402
rect 398932 10338 398984 10344
rect 398944 3398 398972 10338
rect 401324 7812 401376 7818
rect 401324 7754 401376 7760
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 7754
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 39306
rect 405738 17368 405794 17377
rect 405738 17303 405794 17312
rect 405752 16574 405780 17303
rect 408512 16574 408540 62902
rect 412640 61464 412692 61470
rect 412640 61406 412692 61412
rect 411260 43444 411312 43450
rect 411260 43386 411312 43392
rect 411272 16574 411300 43386
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 406028 480 406056 16546
rect 407210 14648 407266 14657
rect 407210 14583 407266 14592
rect 407224 480 407252 14583
rect 408406 8936 408462 8945
rect 408406 8871 408462 8880
rect 408420 480 408448 8871
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 6520 410852 6526
rect 410800 6462 410852 6468
rect 410812 480 410840 6462
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 61406
rect 418160 40724 418212 40730
rect 418160 40666 418212 40672
rect 415400 17604 415452 17610
rect 415400 17546 415452 17552
rect 414296 11892 414348 11898
rect 414296 11834 414348 11840
rect 414308 480 414336 11834
rect 415412 3398 415440 17546
rect 418172 16574 418200 40666
rect 422298 24168 422354 24177
rect 422298 24103 422354 24112
rect 419540 17536 419592 17542
rect 419540 17478 419592 17484
rect 419552 16574 419580 17478
rect 422312 16574 422340 24103
rect 423678 18728 423734 18737
rect 423678 18663 423734 18672
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 417424 13252 417476 13258
rect 417424 13194 417476 13200
rect 415492 11824 415544 11830
rect 415492 11766 415544 11772
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 11766
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 13194
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420918 15872 420974 15881
rect 420918 15807 420974 15816
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15807
rect 422588 480 422616 16546
rect 423692 3210 423720 18663
rect 426452 16574 426480 69838
rect 427820 68400 427872 68406
rect 427820 68342 427872 68348
rect 427832 16574 427860 68342
rect 430592 16574 430620 80038
rect 444380 78804 444432 78810
rect 444380 78746 444432 78752
rect 431960 75540 432012 75546
rect 431960 75482 432012 75488
rect 431972 16574 432000 75482
rect 438860 75472 438912 75478
rect 438860 75414 438912 75420
rect 437480 67108 437532 67114
rect 437480 67050 437532 67056
rect 433340 60036 433392 60042
rect 433340 59978 433392 59984
rect 433352 16574 433380 59978
rect 434720 32700 434772 32706
rect 434720 32642 434772 32648
rect 434732 16574 434760 32642
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 425704 15972 425756 15978
rect 425704 15914 425756 15920
rect 423770 11792 423826 11801
rect 423770 11727 423826 11736
rect 423784 3398 423812 11727
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 15914
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429200 13184 429252 13190
rect 429200 13126 429252 13132
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 13126
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 433248 6452 433300 6458
rect 433248 6394 433300 6400
rect 433260 480 433288 6394
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 14544 436796 14550
rect 436744 14486 436796 14492
rect 436756 480 436784 14486
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 67050
rect 438872 16574 438900 75414
rect 442998 21584 443054 21593
rect 442998 21519 443054 21528
rect 440240 17468 440292 17474
rect 440240 17410 440292 17416
rect 440252 16574 440280 17410
rect 443012 16574 443040 21519
rect 444392 16574 444420 78746
rect 462332 78713 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 142866 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 504364 271924 504416 271930
rect 504364 271866 504416 271872
rect 477500 142860 477552 142866
rect 477500 142802 477552 142808
rect 504376 80889 504404 271866
rect 504456 191888 504508 191894
rect 504456 191830 504508 191836
rect 504362 80880 504418 80889
rect 504362 80815 504418 80824
rect 504468 80714 504496 191830
rect 504456 80708 504508 80714
rect 504456 80650 504508 80656
rect 462318 78704 462374 78713
rect 462318 78639 462374 78648
rect 471980 78124 472032 78130
rect 471980 78066 472032 78072
rect 454040 76560 454092 76566
rect 454040 76502 454092 76508
rect 447140 21616 447192 21622
rect 447140 21558 447192 21564
rect 447152 16574 447180 21558
rect 448520 18896 448572 18902
rect 448520 18838 448572 18844
rect 438872 16546 439176 16574
rect 440252 16546 440372 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 447152 16546 447456 16574
rect 439148 480 439176 16546
rect 440344 480 440372 16546
rect 441528 6384 441580 6390
rect 441528 6326 441580 6332
rect 441540 480 441568 6326
rect 442630 4992 442686 5001
rect 442630 4927 442686 4936
rect 442644 480 442672 4927
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 446220 7744 446272 7750
rect 446220 7686 446272 7692
rect 446232 480 446260 7686
rect 447428 480 447456 16546
rect 448532 3210 448560 18838
rect 451280 18828 451332 18834
rect 451280 18770 451332 18776
rect 448612 17400 448664 17406
rect 448612 17342 448664 17348
rect 448624 3398 448652 17342
rect 451292 16574 451320 18770
rect 451292 16546 451688 16574
rect 450912 5024 450964 5030
rect 450912 4966 450964 4972
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 4966
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453304 13116 453356 13122
rect 453304 13058 453356 13064
rect 453316 480 453344 13058
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 76502
rect 467840 75404 467892 75410
rect 467840 75346 467892 75352
rect 462320 67040 462372 67046
rect 462320 66982 462372 66988
rect 459558 61432 459614 61441
rect 459558 61367 459614 61376
rect 456800 20188 456852 20194
rect 456800 20130 456852 20136
rect 455420 20052 455472 20058
rect 455420 19994 455472 20000
rect 455432 16574 455460 19994
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 20130
rect 458178 20088 458234 20097
rect 458178 20023 458234 20032
rect 456890 17232 456946 17241
rect 456890 17167 456946 17176
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 17167
rect 458192 16574 458220 20023
rect 459572 16574 459600 61367
rect 460938 21448 460994 21457
rect 460938 21383 460994 21392
rect 460952 16574 460980 21383
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 66982
rect 463700 32632 463752 32638
rect 463700 32574 463752 32580
rect 463712 16574 463740 32574
rect 467104 24336 467156 24342
rect 467104 24278 467156 24284
rect 465080 20120 465132 20126
rect 465080 20062 465132 20068
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 6914 465120 20062
rect 465172 19984 465224 19990
rect 465172 19926 465224 19932
rect 465184 16574 465212 19926
rect 465184 16546 465856 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467116 3942 467144 24278
rect 467852 16574 467880 75346
rect 471992 16574 472020 78066
rect 480260 78056 480312 78062
rect 478878 78024 478934 78033
rect 480260 77998 480312 78004
rect 478878 77959 478934 77968
rect 473360 21548 473412 21554
rect 473360 21490 473412 21496
rect 473372 16574 473400 21490
rect 476118 21312 476174 21321
rect 476118 21247 476174 21256
rect 476132 16574 476160 21247
rect 467852 16546 468248 16574
rect 471992 16546 472296 16574
rect 473372 16546 473492 16574
rect 476132 16546 476528 16574
rect 467472 6316 467524 6322
rect 467472 6258 467524 6264
rect 467104 3936 467156 3942
rect 467104 3878 467156 3884
rect 467484 480 467512 6258
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 471060 9104 471112 9110
rect 471060 9046 471112 9052
rect 469864 7676 469916 7682
rect 469864 7618 469916 7624
rect 469876 480 469904 7618
rect 471072 480 471100 9046
rect 472268 480 472296 16546
rect 473464 480 473492 16546
rect 474094 11656 474150 11665
rect 474094 11591 474150 11600
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 11591
rect 475752 3800 475804 3806
rect 475752 3742 475804 3748
rect 475764 480 475792 3742
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478142 14512 478198 14521
rect 478142 14447 478198 14456
rect 478156 480 478184 14447
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 77959
rect 480272 16574 480300 77998
rect 498200 77988 498252 77994
rect 498200 77930 498252 77936
rect 483018 77888 483074 77897
rect 483018 77823 483074 77832
rect 481640 57316 481692 57322
rect 481640 57258 481692 57264
rect 480272 16546 480576 16574
rect 480548 480 480576 16546
rect 481652 6914 481680 57258
rect 481732 32564 481784 32570
rect 481732 32506 481784 32512
rect 481744 16574 481772 32506
rect 483032 16574 483060 77823
rect 490012 75336 490064 75342
rect 490012 75278 490064 75284
rect 496818 75304 496874 75313
rect 488540 62892 488592 62898
rect 488540 62834 488592 62840
rect 484400 21480 484452 21486
rect 484400 21422 484452 21428
rect 484412 16574 484440 21422
rect 488552 16574 488580 62834
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 481652 6886 481772 6914
rect 481744 480 481772 6886
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 10328 486476 10334
rect 486424 10270 486476 10276
rect 486436 480 486464 10270
rect 487620 4956 487672 4962
rect 487620 4898 487672 4904
rect 487632 480 487660 4898
rect 488828 480 488856 16546
rect 490024 6914 490052 75278
rect 496818 75239 496874 75248
rect 494058 71088 494114 71097
rect 494058 71023 494114 71032
rect 492680 17332 492732 17338
rect 492680 17274 492732 17280
rect 492692 16574 492720 17274
rect 494072 16574 494100 71023
rect 495438 19952 495494 19961
rect 495438 19887 495494 19896
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 492312 9036 492364 9042
rect 492312 8978 492364 8984
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3732 491168 3738
rect 491116 3674 491168 3680
rect 491128 480 491156 3674
rect 492324 480 492352 8978
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 19887
rect 496832 16574 496860 75239
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 77930
rect 527192 77246 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 141574 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 579986 458144 580042 458153
rect 579986 458079 580042 458088
rect 580000 456822 580028 458079
rect 579988 456816 580040 456822
rect 579988 456758 580040 456764
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580092 418198 580120 418231
rect 580080 418192 580132 418198
rect 580080 418134 580132 418140
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580092 378214 580120 378383
rect 580080 378208 580132 378214
rect 580080 378150 580132 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580092 311914 580120 312015
rect 580080 311908 580132 311914
rect 580080 311850 580132 311856
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580092 298178 580120 298687
rect 580080 298172 580132 298178
rect 580080 298114 580132 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 580092 231878 580120 232319
rect 580080 231872 580132 231878
rect 580080 231814 580132 231820
rect 580078 219056 580134 219065
rect 580078 218991 580134 219000
rect 580092 218074 580120 218991
rect 580080 218068 580132 218074
rect 580080 218010 580132 218016
rect 580078 205728 580134 205737
rect 580078 205663 580080 205672
rect 580132 205663 580134 205672
rect 580080 205634 580132 205640
rect 579802 192536 579858 192545
rect 579802 192471 579858 192480
rect 579816 191894 579844 192471
rect 579804 191888 579856 191894
rect 579804 191830 579856 191836
rect 580078 179208 580134 179217
rect 580078 179143 580134 179152
rect 580092 175982 580120 179143
rect 580080 175976 580132 175982
rect 580080 175918 580132 175924
rect 580078 165880 580134 165889
rect 580078 165815 580134 165824
rect 580092 165646 580120 165815
rect 580080 165640 580132 165646
rect 580080 165582 580132 165588
rect 580184 158030 580212 471407
rect 580172 158024 580224 158030
rect 580172 157966 580224 157972
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 542360 141568 542412 141574
rect 542360 141510 542412 141516
rect 580276 141506 580304 683839
rect 580722 630864 580778 630873
rect 580722 630799 580778 630808
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 141500 580316 141506
rect 580264 141442 580316 141448
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580184 125662 580212 125967
rect 580172 125656 580224 125662
rect 580172 125598 580224 125604
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 555424 81456 555476 81462
rect 580276 81433 580304 99447
rect 580368 82142 580396 590951
rect 580538 577688 580594 577697
rect 580538 577623 580594 577632
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580356 82136 580408 82142
rect 580356 82078 580408 82084
rect 555424 81398 555476 81404
rect 580262 81424 580318 81433
rect 554780 78736 554832 78742
rect 554780 78678 554832 78684
rect 527180 77240 527232 77246
rect 527180 77182 527232 77188
rect 549258 76664 549314 76673
rect 549258 76599 549314 76608
rect 499580 75268 499632 75274
rect 499580 75210 499632 75216
rect 498292 23112 498344 23118
rect 498292 23054 498344 23060
rect 498304 16574 498332 23054
rect 499592 16574 499620 75210
rect 528558 75168 528614 75177
rect 528558 75103 528614 75112
rect 505100 69828 505152 69834
rect 505100 69770 505152 69776
rect 505112 16574 505140 69770
rect 518900 69760 518952 69766
rect 518900 69702 518952 69708
rect 511998 68232 512054 68241
rect 511998 68167 512054 68176
rect 507860 57248 507912 57254
rect 507860 57190 507912 57196
rect 506480 26920 506532 26926
rect 506480 26862 506532 26868
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 505112 16546 505416 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 502984 14476 503036 14482
rect 502984 14418 503036 14424
rect 501788 3664 501840 3670
rect 501788 3606 501840 3612
rect 501800 480 501828 3606
rect 502996 480 503024 14418
rect 504180 7608 504232 7614
rect 504180 7550 504232 7556
rect 504192 480 504220 7550
rect 505388 480 505416 16546
rect 506492 3398 506520 26862
rect 506572 21412 506624 21418
rect 506572 21354 506624 21360
rect 506480 3392 506532 3398
rect 506480 3334 506532 3340
rect 506584 3210 506612 21354
rect 507872 16574 507900 57190
rect 510618 27024 510674 27033
rect 510618 26959 510674 26968
rect 509240 23044 509292 23050
rect 509240 22986 509292 22992
rect 509252 16574 509280 22986
rect 510632 16574 510660 26959
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511304 16574
rect 507308 3392 507360 3398
rect 507308 3334 507360 3340
rect 506492 3182 506612 3210
rect 506492 480 506520 3182
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3334
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511276 480 511304 16546
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 68167
rect 514850 28248 514906 28257
rect 514850 28183 514906 28192
rect 513378 10296 513434 10305
rect 513378 10231 513434 10240
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 10231
rect 514864 6914 514892 28183
rect 517520 25764 517572 25770
rect 517520 25706 517572 25712
rect 516140 22976 516192 22982
rect 516140 22918 516192 22924
rect 516152 16574 516180 22918
rect 517532 16574 517560 25706
rect 518912 16574 518940 69702
rect 525800 61396 525852 61402
rect 525800 61338 525852 61344
rect 524420 31068 524472 31074
rect 524420 31010 524472 31016
rect 521660 29708 521712 29714
rect 521660 29650 521712 29656
rect 520280 22908 520332 22914
rect 520280 22850 520332 22856
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 514772 6886 514892 6914
rect 514772 480 514800 6886
rect 515956 3596 516008 3602
rect 515956 3538 516008 3544
rect 515968 480 515996 3538
rect 517164 480 517192 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22850
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 29650
rect 524432 16574 524460 31010
rect 525812 16574 525840 61338
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523776 11756 523828 11762
rect 523776 11698 523828 11704
rect 523040 4888 523092 4894
rect 523040 4830 523092 4836
rect 523052 480 523080 4830
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 11698
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 4820 527876 4826
rect 527824 4762 527876 4768
rect 527836 480 527864 4762
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 75103
rect 539600 66972 539652 66978
rect 539600 66914 539652 66920
rect 529938 62928 529994 62937
rect 529938 62863 529994 62872
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 62863
rect 531318 32600 531374 32609
rect 531318 32535 531374 32544
rect 531332 3534 531360 32535
rect 535460 24268 535512 24274
rect 535460 24210 535512 24216
rect 535472 16574 535500 24210
rect 538220 24200 538272 24206
rect 538220 24142 538272 24148
rect 535472 16546 536144 16574
rect 531410 13016 531466 13025
rect 531410 12951 531466 12960
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 12951
rect 534908 3936 534960 3942
rect 534908 3878 534960 3884
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 534920 480 534948 3878
rect 536116 480 536144 16546
rect 537208 3392 537260 3398
rect 537208 3334 537260 3340
rect 537220 480 537248 3334
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24142
rect 539612 3534 539640 66914
rect 543740 66904 543792 66910
rect 543740 66846 543792 66852
rect 539692 32496 539744 32502
rect 539692 32438 539744 32444
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 32438
rect 542360 29640 542412 29646
rect 542360 29582 542412 29588
rect 542372 16574 542400 29582
rect 543752 16574 543780 66846
rect 546498 30968 546554 30977
rect 546498 30903 546554 30912
rect 545120 17264 545172 17270
rect 545120 17206 545172 17212
rect 545132 16574 545160 17206
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 541992 15904 542044 15910
rect 541992 15846 542044 15852
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 15846
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 30903
rect 547878 18592 547934 18601
rect 547878 18527 547934 18536
rect 547892 16574 547920 18527
rect 549272 16574 549300 76599
rect 550638 62792 550694 62801
rect 550638 62727 550694 62736
rect 550652 16574 550680 62727
rect 552020 24132 552072 24138
rect 552020 24074 552072 24080
rect 552032 16574 552060 24074
rect 553400 18760 553452 18766
rect 553400 18702 553452 18708
rect 553412 16574 553440 18702
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 547878 4856 547934 4865
rect 547878 4791 547934 4800
rect 547892 480 547920 4791
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 78678
rect 555436 6866 555464 81398
rect 580262 81359 580318 81368
rect 580460 79354 580488 537775
rect 580552 141438 580580 577623
rect 580630 484664 580686 484673
rect 580630 484599 580686 484608
rect 580540 141432 580592 141438
rect 580540 141374 580592 141380
rect 580448 79348 580500 79354
rect 580448 79290 580500 79296
rect 580644 77586 580672 484599
rect 580736 228410 580764 630799
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580724 228404 580776 228410
rect 580724 228346 580776 228352
rect 580828 164898 580856 524447
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580816 164892 580868 164898
rect 580816 164834 580868 164840
rect 580920 80753 580948 431559
rect 580906 80744 580962 80753
rect 580906 80679 580962 80688
rect 580632 77580 580684 77586
rect 580632 77522 580684 77528
rect 565818 76528 565874 76537
rect 565818 76463 565874 76472
rect 564440 75200 564492 75206
rect 564440 75142 564492 75148
rect 561680 64184 561732 64190
rect 561680 64126 561732 64132
rect 557540 62824 557592 62830
rect 557540 62766 557592 62772
rect 556160 22840 556212 22846
rect 556160 22782 556212 22788
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 556172 480 556200 22782
rect 556252 18692 556304 18698
rect 556252 18634 556304 18640
rect 556264 16574 556292 18634
rect 557552 16574 557580 62766
rect 558920 25696 558972 25702
rect 558920 25638 558972 25644
rect 558932 16574 558960 25638
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 561692 16574 561720 64126
rect 563060 25628 563112 25634
rect 563060 25570 563112 25576
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 25570
rect 564452 480 564480 75142
rect 564532 68332 564584 68338
rect 564532 68274 564584 68280
rect 564544 16574 564572 68274
rect 565832 16574 565860 76463
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 568580 69692 568632 69698
rect 568580 69634 568632 69640
rect 567198 32464 567254 32473
rect 567198 32399 567254 32408
rect 567212 16574 567240 32399
rect 568592 16574 568620 69634
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 578238 33824 578294 33833
rect 578238 33759 578294 33768
rect 574100 32428 574152 32434
rect 574100 32370 574152 32376
rect 572720 25560 572772 25566
rect 572720 25502 572772 25508
rect 572732 16574 572760 25502
rect 574112 16574 574140 32370
rect 576858 26888 576914 26897
rect 576858 26823 576914 26832
rect 576872 16574 576900 26823
rect 578252 16574 578280 33759
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 581000 28280 581052 28286
rect 581000 28222 581052 28228
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 581012 16574 581040 28222
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 572732 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 581012 16546 581776 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 571524 8968 571576 8974
rect 571524 8910 571576 8916
rect 570326 3496 570382 3505
rect 570326 3431 570382 3440
rect 570340 480 570368 3431
rect 571536 480 571564 8910
rect 572720 6248 572772 6254
rect 572720 6190 572772 6196
rect 572732 480 572760 6190
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 576320 480 576348 6122
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 3868 583444 3874
rect 583392 3810 583444 3816
rect 583404 480 583432 3810
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3054 566888 3110 566944
rect 2962 527856 3018 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3330 423544 3386 423600
rect 3238 410508 3294 410544
rect 3238 410488 3240 410508
rect 3240 410488 3292 410508
rect 3292 410488 3294 410508
rect 3238 371320 3294 371376
rect 3238 358400 3294 358456
rect 3238 319232 3294 319288
rect 3238 306176 3294 306232
rect 2778 293120 2834 293176
rect 3054 267144 3110 267200
rect 3146 254088 3202 254144
rect 2778 241032 2834 241088
rect 2870 227976 2926 228032
rect 3330 214920 3386 214976
rect 3330 201884 3386 201920
rect 3330 201864 3332 201884
rect 3332 201864 3384 201884
rect 3384 201864 3386 201884
rect 3330 188808 3386 188864
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 3330 136720 3386 136776
rect 3146 110608 3202 110664
rect 3238 97552 3294 97608
rect 3514 619112 3570 619168
rect 3606 606056 3662 606112
rect 3514 579944 3570 580000
rect 3514 553832 3570 553888
rect 3790 501744 3846 501800
rect 3698 449520 3754 449576
rect 3146 80416 3202 80472
rect 3238 78920 3294 78976
rect 1398 76472 1454 76528
rect 2778 75112 2834 75168
rect 3514 81232 3570 81288
rect 4066 475632 4122 475688
rect 3974 397432 4030 397488
rect 3882 345344 3938 345400
rect 4066 149776 4122 149832
rect 3974 84632 4030 84688
rect 3882 80552 3938 80608
rect 3790 79328 3846 79384
rect 3606 79192 3662 79248
rect 3422 79056 3478 79112
rect 3422 71576 3478 71632
rect 3330 58520 3386 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 6918 79464 6974 79520
rect 117318 136856 117374 136912
rect 117318 135360 117374 135416
rect 117318 133900 117320 133920
rect 117320 133900 117372 133920
rect 117372 133900 117374 133920
rect 117318 133864 117374 133900
rect 117318 132404 117320 132424
rect 117320 132404 117372 132424
rect 117372 132404 117374 132424
rect 117318 132368 117374 132404
rect 117318 130872 117374 130928
rect 117318 129376 117374 129432
rect 117318 127880 117374 127936
rect 117318 126384 117374 126440
rect 117318 124888 117374 124944
rect 117318 123392 117374 123448
rect 117318 121896 117374 121952
rect 117318 120400 117374 120456
rect 117318 118904 117374 118960
rect 117318 117408 117374 117464
rect 117318 115912 117374 115968
rect 117318 114452 117320 114472
rect 117320 114452 117372 114472
rect 117372 114452 117374 114472
rect 117318 114416 117374 114452
rect 117318 112920 117374 112976
rect 117318 111424 117374 111480
rect 117318 109928 117374 109984
rect 118054 108432 118110 108488
rect 117870 106936 117926 106992
rect 118146 103944 118202 104000
rect 118238 94968 118294 95024
rect 118330 93472 118386 93528
rect 118422 91976 118478 92032
rect 118514 90480 118570 90536
rect 138110 195916 138112 195936
rect 138112 195916 138164 195936
rect 138164 195916 138166 195936
rect 138110 195880 138166 195916
rect 140410 195880 140466 195936
rect 158810 195872 158866 195928
rect 160098 195916 160100 195936
rect 160100 195916 160152 195936
rect 160152 195916 160154 195936
rect 160098 195880 160154 195916
rect 140778 195608 140834 195664
rect 139398 195472 139454 195528
rect 140870 191800 140926 191856
rect 140778 191528 140834 191584
rect 140962 190848 141018 190904
rect 140870 184320 140926 184376
rect 140778 184184 140834 184240
rect 140962 184048 141018 184104
rect 118790 100952 118846 101008
rect 118698 88984 118754 89040
rect 118974 97960 119030 98016
rect 119250 102448 119306 102504
rect 119158 99456 119214 99512
rect 119066 96464 119122 96520
rect 118882 87488 118938 87544
rect 118606 85992 118662 86048
rect 118514 83000 118570 83056
rect 118422 81504 118478 81560
rect 20718 76608 20774 76664
rect 4066 19352 4122 19408
rect 22098 43424 22154 43480
rect 3422 6432 3478 6488
rect 4066 4800 4122 4856
rect 20626 3304 20682 3360
rect 35898 75248 35954 75304
rect 40038 73752 40094 73808
rect 38382 7520 38438 7576
rect 41878 7656 41934 7712
rect 53838 75384 53894 75440
rect 57150 8880 57206 8936
rect 56046 7792 56102 7848
rect 57978 75520 58034 75576
rect 111798 76880 111854 76936
rect 93858 76744 93914 76800
rect 91098 44784 91154 44840
rect 73802 6160 73858 6216
rect 72606 3440 72662 3496
rect 78586 9016 78642 9072
rect 92478 10240 92534 10296
rect 144366 190984 144422 191040
rect 145838 188944 145894 189000
rect 144918 188128 144974 188184
rect 144918 181192 144974 181248
rect 144642 180920 144698 180976
rect 157798 179444 157854 179480
rect 157798 179424 157800 179444
rect 157800 179424 157852 179444
rect 157852 179424 157854 179444
rect 158534 179424 158590 179480
rect 144090 178880 144146 178936
rect 143078 178744 143134 178800
rect 141606 178608 141662 178664
rect 163502 175888 163558 175944
rect 149334 175616 149390 175672
rect 158166 175616 158222 175672
rect 165158 175908 165214 175944
rect 165158 175888 165160 175908
rect 165160 175888 165212 175908
rect 165212 175888 165214 175908
rect 163594 175752 163650 175808
rect 165066 175752 165122 175808
rect 155222 171808 155278 171864
rect 171506 142840 171562 142896
rect 173070 142704 173126 142760
rect 121274 138896 121330 138952
rect 179602 135496 179658 135552
rect 179510 131960 179566 132016
rect 179418 126112 179474 126168
rect 120630 105984 120686 106040
rect 120630 84224 120686 84280
rect 120630 81368 120686 81424
rect 110510 10376 110566 10432
rect 109314 7928 109370 7984
rect 111614 6296 111670 6352
rect 178406 80960 178462 81016
rect 178314 80824 178370 80880
rect 123022 79736 123078 79792
rect 123666 75248 123722 75304
rect 174634 80300 174690 80336
rect 174634 80280 174636 80300
rect 174636 80280 174688 80300
rect 174688 80280 174690 80300
rect 125736 79872 125792 79928
rect 126104 79872 126160 79928
rect 126380 79906 126436 79962
rect 127116 79906 127172 79962
rect 125690 76472 125746 76528
rect 125782 75928 125838 75984
rect 126150 79600 126206 79656
rect 127300 79872 127356 79928
rect 127852 79906 127908 79962
rect 127714 79736 127770 79792
rect 128128 79906 128184 79962
rect 127070 44920 127126 44976
rect 127254 76608 127310 76664
rect 127530 79600 127586 79656
rect 127990 78104 128046 78160
rect 128496 79906 128552 79962
rect 128680 79906 128736 79962
rect 128864 79906 128920 79962
rect 129232 79872 129288 79928
rect 130060 79872 130116 79928
rect 130336 79872 130392 79928
rect 128358 76472 128414 76528
rect 128726 77968 128782 78024
rect 127990 73752 128046 73808
rect 129186 79600 129242 79656
rect 129738 77968 129794 78024
rect 130014 78104 130070 78160
rect 130106 77968 130162 78024
rect 130474 77968 130530 78024
rect 131256 79906 131312 79962
rect 131440 79906 131496 79962
rect 131624 79906 131680 79962
rect 131900 79906 131956 79962
rect 131394 79736 131450 79792
rect 131026 77968 131082 78024
rect 130382 74432 130438 74488
rect 131854 79600 131910 79656
rect 132360 79906 132416 79962
rect 132636 79906 132692 79962
rect 132314 79736 132370 79792
rect 132498 79600 132554 79656
rect 132866 77424 132922 77480
rect 132590 76744 132646 76800
rect 133464 79838 133520 79894
rect 133832 79872 133888 79928
rect 134200 79906 134256 79962
rect 134384 79906 134440 79962
rect 133786 79600 133842 79656
rect 134016 79736 134072 79792
rect 134338 79736 134394 79792
rect 134844 79872 134900 79928
rect 134062 79636 134064 79656
rect 134064 79636 134116 79656
rect 134116 79636 134118 79656
rect 134062 79600 134118 79636
rect 134154 76880 134210 76936
rect 134798 79736 134854 79792
rect 135396 79872 135452 79928
rect 135764 79872 135820 79928
rect 135718 79736 135774 79792
rect 135534 77968 135590 78024
rect 136040 79906 136096 79962
rect 137144 79906 137200 79962
rect 137328 79906 137384 79962
rect 136086 79600 136142 79656
rect 137190 79736 137246 79792
rect 137558 79736 137614 79792
rect 137972 79736 138028 79792
rect 138432 79906 138488 79962
rect 138984 79872 139040 79928
rect 139536 79872 139592 79928
rect 137834 78104 137890 78160
rect 138018 77968 138074 78024
rect 138570 78784 138626 78840
rect 139168 79736 139224 79792
rect 139582 79736 139638 79792
rect 139996 79906 140052 79962
rect 139398 79600 139454 79656
rect 139122 75656 139178 75712
rect 139950 79756 140006 79792
rect 139950 79736 139952 79756
rect 139952 79736 140004 79756
rect 140004 79736 140006 79756
rect 140640 79872 140696 79928
rect 141100 79906 141156 79962
rect 139950 79600 140006 79656
rect 139950 75520 140006 75576
rect 140410 75792 140466 75848
rect 140594 75928 140650 75984
rect 142020 79906 142076 79962
rect 140686 74024 140742 74080
rect 142756 79906 142812 79962
rect 142526 79736 142582 79792
rect 143308 79906 143364 79962
rect 142066 79600 142122 79656
rect 142618 76064 142674 76120
rect 142848 79736 142904 79792
rect 143492 79872 143548 79928
rect 142894 79600 142950 79656
rect 143262 79636 143264 79656
rect 143264 79636 143316 79656
rect 143316 79636 143318 79656
rect 143262 79600 143318 79636
rect 143952 79906 144008 79962
rect 144320 79872 144376 79928
rect 144596 79872 144652 79928
rect 144872 79906 144928 79962
rect 145056 79838 145112 79894
rect 143262 75928 143318 75984
rect 143722 79600 143778 79656
rect 143814 75928 143870 75984
rect 144642 78648 144698 78704
rect 144734 76880 144790 76936
rect 145102 79600 145158 79656
rect 145516 79872 145572 79928
rect 145976 79872 146032 79928
rect 145470 79600 145526 79656
rect 146160 79872 146216 79928
rect 145930 78784 145986 78840
rect 146344 79872 146400 79928
rect 146206 78648 146262 78704
rect 146114 78512 146170 78568
rect 147356 79906 147412 79962
rect 148000 79872 148056 79928
rect 147632 79770 147688 79826
rect 147402 78648 147458 78704
rect 147678 76744 147734 76800
rect 148736 79872 148792 79928
rect 148920 79736 148976 79792
rect 148966 79600 149022 79656
rect 148782 78648 148838 78704
rect 149058 78784 149114 78840
rect 149058 78648 149114 78704
rect 148874 78376 148930 78432
rect 148874 77424 148930 77480
rect 149840 79872 149896 79928
rect 150208 79838 150264 79894
rect 150392 79838 150448 79894
rect 151036 79872 151092 79928
rect 149702 78784 149758 78840
rect 150254 78648 150310 78704
rect 150438 78648 150494 78704
rect 150162 78512 150218 78568
rect 150852 79736 150908 79792
rect 151312 79906 151368 79962
rect 151772 79872 151828 79928
rect 152232 79906 152288 79962
rect 151726 79736 151782 79792
rect 150990 77832 151046 77888
rect 152186 79736 152242 79792
rect 152416 79906 152472 79962
rect 152600 79872 152656 79928
rect 151174 78648 151230 78704
rect 151358 78784 151414 78840
rect 151726 78512 151782 78568
rect 152002 79600 152058 79656
rect 152646 79736 152702 79792
rect 152876 79872 152932 79928
rect 153152 79906 153208 79962
rect 153014 79736 153070 79792
rect 152830 76608 152886 76664
rect 153106 79600 153162 79656
rect 153014 77288 153070 77344
rect 153888 79906 153944 79962
rect 154440 79906 154496 79962
rect 154210 78648 154266 78704
rect 154394 75928 154450 75984
rect 154670 79736 154726 79792
rect 154900 79872 154956 79928
rect 155084 79906 155140 79962
rect 155544 79906 155600 79962
rect 154486 75792 154542 75848
rect 155038 79736 155094 79792
rect 155728 79872 155784 79928
rect 156096 79872 156152 79928
rect 155866 79736 155922 79792
rect 156648 79872 156704 79928
rect 157108 79872 157164 79928
rect 157292 79906 157348 79962
rect 155038 78104 155094 78160
rect 155222 75928 155278 75984
rect 155682 79600 155738 79656
rect 155866 76200 155922 76256
rect 156372 79736 156428 79792
rect 156050 79600 156106 79656
rect 156142 75928 156198 75984
rect 156418 77832 156474 77888
rect 156786 79600 156842 79656
rect 156878 75384 156934 75440
rect 157246 78784 157302 78840
rect 157154 78240 157210 78296
rect 157062 77424 157118 77480
rect 158396 79872 158452 79928
rect 158580 79872 158636 79928
rect 158948 79906 159004 79962
rect 159776 79906 159832 79962
rect 158534 78104 158590 78160
rect 158442 77968 158498 78024
rect 158810 78512 158866 78568
rect 159178 77968 159234 78024
rect 160052 79906 160108 79962
rect 160512 79906 160568 79962
rect 159730 78648 159786 78704
rect 160282 78648 160338 78704
rect 160880 79906 160936 79962
rect 161340 79906 161396 79962
rect 161524 79906 161580 79962
rect 161294 79736 161350 79792
rect 161984 79872 162040 79928
rect 160926 79600 160982 79656
rect 161018 78648 161074 78704
rect 161386 79600 161442 79656
rect 161202 78512 161258 78568
rect 161202 77968 161258 78024
rect 161570 78648 161626 78704
rect 161478 78376 161534 78432
rect 160558 19896 160614 19952
rect 158902 4800 158958 4856
rect 161846 79600 161902 79656
rect 162398 79736 162454 79792
rect 162628 79872 162684 79928
rect 162720 79736 162776 79792
rect 162996 79906 163052 79962
rect 162122 78376 162178 78432
rect 162490 78648 162546 78704
rect 162214 77152 162270 77208
rect 162674 78648 162730 78704
rect 162950 79736 163006 79792
rect 163180 79906 163236 79962
rect 163548 79906 163604 79962
rect 163824 79872 163880 79928
rect 164008 79906 164064 79962
rect 162858 77968 162914 78024
rect 161294 3304 161350 3360
rect 163364 79736 163420 79792
rect 163226 78648 163282 78704
rect 163134 77560 163190 77616
rect 163870 79736 163926 79792
rect 164284 79872 164340 79928
rect 163502 78784 163558 78840
rect 163594 77696 163650 77752
rect 164560 79906 164616 79962
rect 164238 79600 164294 79656
rect 164146 75248 164202 75304
rect 165296 79906 165352 79962
rect 164790 78648 164846 78704
rect 165066 77560 165122 77616
rect 165572 79906 165628 79962
rect 165342 79600 165398 79656
rect 165434 78784 165490 78840
rect 165710 79620 165766 79656
rect 165710 79600 165712 79620
rect 165712 79600 165764 79620
rect 165764 79600 165766 79620
rect 165618 78648 165674 78704
rect 165526 78512 165582 78568
rect 165802 78648 165858 78704
rect 166216 79736 166272 79792
rect 166400 79736 166456 79792
rect 166262 79600 166318 79656
rect 166676 79872 166732 79928
rect 167320 79872 167376 79928
rect 166722 78648 166778 78704
rect 166630 78104 166686 78160
rect 166630 77696 166686 77752
rect 166906 79620 166962 79656
rect 166906 79600 166908 79620
rect 166908 79600 166960 79620
rect 166960 79600 166962 79620
rect 166814 77560 166870 77616
rect 167090 78104 167146 78160
rect 167688 79872 167744 79928
rect 167872 79872 167928 79928
rect 167642 78512 167698 78568
rect 168240 79872 168296 79928
rect 168424 79872 168480 79928
rect 168792 79906 168848 79962
rect 168976 79872 169032 79928
rect 168562 79736 168618 79792
rect 168838 79736 168894 79792
rect 169022 79736 169078 79792
rect 168010 78648 168066 78704
rect 168194 78104 168250 78160
rect 168102 77560 168158 77616
rect 168746 78376 168802 78432
rect 168654 78104 168710 78160
rect 168930 78104 168986 78160
rect 168838 76472 168894 76528
rect 169436 79872 169492 79928
rect 169620 79872 169676 79928
rect 169574 78512 169630 78568
rect 169896 79906 169952 79962
rect 170080 79906 170136 79962
rect 170264 79872 170320 79928
rect 170448 79872 170504 79928
rect 169666 78104 169722 78160
rect 169850 78648 169906 78704
rect 170724 79872 170780 79928
rect 170908 79872 170964 79928
rect 170126 79600 170182 79656
rect 170310 79600 170366 79656
rect 170494 79600 170550 79656
rect 170218 78104 170274 78160
rect 170218 77832 170274 77888
rect 171184 79872 171240 79928
rect 171460 79906 171516 79962
rect 171644 79872 171700 79928
rect 170218 77016 170274 77072
rect 170218 76608 170274 76664
rect 170586 78648 170642 78704
rect 170862 78668 170918 78704
rect 170862 78648 170864 78668
rect 170864 78648 170916 78668
rect 170916 78648 170918 78668
rect 170862 78512 170918 78568
rect 171046 79600 171102 79656
rect 171598 79736 171654 79792
rect 171506 79600 171562 79656
rect 172288 79872 172344 79928
rect 172472 79872 172528 79928
rect 171506 78376 171562 78432
rect 171138 75928 171194 75984
rect 171782 78668 171838 78704
rect 171782 78648 171784 78668
rect 171784 78648 171836 78668
rect 171836 78648 171838 78668
rect 172150 78648 172206 78704
rect 172748 79736 172804 79792
rect 172334 78648 172390 78704
rect 172242 78512 172298 78568
rect 171966 77288 172022 77344
rect 171874 77172 171930 77208
rect 171874 77152 171876 77172
rect 171876 77152 171928 77172
rect 171928 77152 171930 77172
rect 172334 78240 172390 78296
rect 172242 78104 172298 78160
rect 172702 78376 172758 78432
rect 173300 79872 173356 79928
rect 172978 79464 173034 79520
rect 173760 79872 173816 79928
rect 173346 79192 173402 79248
rect 173668 79772 173670 79792
rect 173670 79772 173722 79792
rect 173722 79772 173724 79792
rect 173668 79736 173724 79772
rect 173254 79056 173310 79112
rect 173530 79056 173586 79112
rect 173070 78920 173126 78976
rect 172518 60016 172574 60072
rect 174266 79736 174322 79792
rect 173990 78240 174046 78296
rect 173254 76608 173310 76664
rect 173898 75656 173954 75712
rect 174542 79328 174598 79384
rect 178314 80144 178370 80200
rect 178498 79600 178554 79656
rect 175278 69536 175334 69592
rect 176658 75520 176714 75576
rect 178774 77288 178830 77344
rect 178682 72664 178738 72720
rect 180890 137536 180946 137592
rect 180798 124072 180854 124128
rect 180062 81232 180118 81288
rect 180982 116592 181038 116648
rect 182178 134544 182234 134600
rect 181258 133048 181314 133104
rect 181166 115096 181222 115152
rect 182270 122576 182326 122632
rect 182638 128560 182694 128616
rect 182546 127064 182602 127120
rect 182914 130056 182970 130112
rect 182730 121080 182786 121136
rect 182454 119584 182510 119640
rect 182362 118088 182418 118144
rect 182178 113600 182234 113656
rect 181074 112104 181130 112160
rect 183282 110608 183338 110664
rect 183466 109112 183522 109168
rect 183374 107616 183430 107672
rect 183466 106120 183522 106176
rect 183466 104624 183522 104680
rect 183466 103128 183522 103184
rect 183466 101632 183522 101688
rect 183466 100136 183522 100192
rect 183466 98640 183522 98696
rect 183466 97144 183522 97200
rect 183190 95648 183246 95704
rect 183282 94152 183338 94208
rect 183282 92656 183338 92712
rect 183466 91160 183522 91216
rect 183466 89684 183522 89720
rect 183466 89664 183468 89684
rect 183468 89664 183520 89684
rect 183520 89664 183522 89684
rect 183466 88204 183468 88224
rect 183468 88204 183520 88224
rect 183520 88204 183522 88224
rect 183466 88168 183522 88204
rect 182822 86672 182878 86728
rect 183466 85176 183522 85232
rect 182822 83680 182878 83736
rect 183466 82184 183522 82240
rect 194598 74024 194654 74080
rect 193218 65456 193274 65512
rect 191838 18944 191894 19000
rect 193310 28464 193366 28520
rect 213366 10648 213422 10704
rect 230478 73888 230534 73944
rect 227718 59880 227774 59936
rect 226430 34040 226486 34096
rect 229098 28328 229154 28384
rect 247038 76880 247094 76936
rect 244278 73752 244334 73808
rect 248418 20168 248474 20224
rect 246394 7656 246450 7712
rect 266358 33904 266414 33960
rect 264150 9152 264206 9208
rect 265346 7520 265402 7576
rect 396814 81096 396870 81152
rect 396998 80960 397054 81016
rect 397458 78784 397514 78840
rect 396722 78512 396778 78568
rect 282918 76744 282974 76800
rect 280158 44784 280214 44840
rect 284298 72528 284354 72584
rect 281538 10512 281594 10568
rect 298098 72392 298154 72448
rect 301502 13232 301558 13288
rect 299662 10376 299718 10432
rect 300766 9016 300822 9072
rect 316038 53080 316094 53136
rect 315026 5072 315082 5128
rect 317418 29552 317474 29608
rect 319442 21664 319498 21720
rect 316222 16224 316278 16280
rect 336278 6432 336334 6488
rect 333886 6160 333942 6216
rect 335082 3576 335138 3632
rect 337474 6296 337530 6352
rect 353298 71168 353354 71224
rect 351918 47504 351974 47560
rect 350538 18808 350594 18864
rect 349250 13096 349306 13152
rect 367098 40568 367154 40624
rect 372618 35128 372674 35184
rect 371238 16088 371294 16144
rect 370134 14728 370190 14784
rect 386418 25472 386474 25528
rect 387798 15952 387854 16008
rect 402978 75384 403034 75440
rect 405738 17312 405794 17368
rect 407210 14592 407266 14648
rect 408406 8880 408462 8936
rect 422298 24112 422354 24168
rect 423678 18672 423734 18728
rect 420918 15816 420974 15872
rect 423770 11736 423826 11792
rect 442998 21528 443054 21584
rect 504362 80824 504418 80880
rect 462318 78648 462374 78704
rect 442630 4936 442686 4992
rect 459558 61376 459614 61432
rect 458178 20032 458234 20088
rect 456890 17176 456946 17232
rect 460938 21392 460994 21448
rect 478878 77968 478934 78024
rect 476118 21256 476174 21312
rect 474094 11600 474150 11656
rect 478142 14456 478198 14512
rect 483018 77832 483074 77888
rect 496818 75248 496874 75304
rect 494058 71032 494114 71088
rect 495438 19896 495494 19952
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 617480 580226 617536
rect 580170 564304 580226 564360
rect 580170 511264 580226 511320
rect 580170 471416 580226 471472
rect 579986 458088 580042 458144
rect 580078 418240 580134 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 579802 365064 579858 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 325216 580134 325272
rect 580078 312024 580134 312080
rect 580078 298696 580134 298752
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 580078 232328 580134 232384
rect 580078 219000 580134 219056
rect 580078 205692 580134 205728
rect 580078 205672 580080 205692
rect 580080 205672 580132 205692
rect 580132 205672 580134 205692
rect 579802 192480 579858 192536
rect 580078 179152 580134 179208
rect 580078 165824 580134 165880
rect 579986 152632 580042 152688
rect 580722 630808 580778 630864
rect 580354 590960 580410 591016
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580538 577632 580594 577688
rect 580446 537784 580502 537840
rect 549258 76608 549314 76664
rect 528558 75112 528614 75168
rect 511998 68176 512054 68232
rect 510618 26968 510674 27024
rect 514850 28192 514906 28248
rect 513378 10240 513434 10296
rect 529938 62872 529994 62928
rect 531318 32544 531374 32600
rect 531410 12960 531466 13016
rect 546498 30912 546554 30968
rect 547878 18536 547934 18592
rect 550638 62736 550694 62792
rect 547878 4800 547934 4856
rect 580262 81368 580318 81424
rect 580630 484608 580686 484664
rect 580814 524456 580870 524512
rect 580906 431568 580962 431624
rect 580906 80688 580962 80744
rect 565818 76472 565874 76528
rect 580170 72936 580226 72992
rect 567198 32408 567254 32464
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 578238 33768 578294 33824
rect 576858 26832 576914 26888
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 570326 3440 570382 3496
rect 580170 6568 580226 6624
rect 580998 3304 581054 3360
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 567150 697174 584960 697234
rect 396574 696900 396580 696964
rect 396644 696962 396650 696964
rect 567150 696962 567210 697174
rect 583520 697084 584960 697174
rect 396644 696902 567210 696962
rect 396644 696900 396650 696902
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580717 630866 580783 630869
rect 583520 630866 584960 630956
rect 580717 630864 584960 630866
rect 580717 630808 580722 630864
rect 580778 630808 584960 630864
rect 580717 630806 584960 630808
rect 580717 630803 580783 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580533 577690 580599 577693
rect 583520 577690 584960 577780
rect 580533 577688 584960 577690
rect 580533 577632 580538 577688
rect 580594 577632 584960 577688
rect 580533 577630 584960 577632
rect 580533 577627 580599 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580625 484666 580691 484669
rect 583520 484666 584960 484756
rect 580625 484664 584960 484666
rect 580625 484608 580630 484664
rect 580686 484608 584960 484664
rect 580625 484606 584960 484608
rect 580625 484603 580691 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 4061 475690 4127 475693
rect -960 475688 4127 475690
rect -960 475632 4066 475688
rect 4122 475632 4127 475688
rect -960 475630 4127 475632
rect -960 475540 480 475630
rect 4061 475627 4127 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 579981 458146 580047 458149
rect 583520 458146 584960 458236
rect 579981 458144 584960 458146
rect 579981 458088 579986 458144
rect 580042 458088 584960 458144
rect 579981 458086 584960 458088
rect 579981 458083 580047 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3233 358458 3299 358461
rect -960 358456 3299 358458
rect -960 358400 3238 358456
rect 3294 358400 3299 358456
rect -960 358398 3299 358400
rect -960 358308 480 358398
rect 3233 358395 3299 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3877 345402 3943 345405
rect -960 345400 3943 345402
rect -960 345344 3882 345400
rect 3938 345344 3943 345400
rect -960 345342 3943 345344
rect -960 345252 480 345342
rect 3877 345339 3943 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3233 319290 3299 319293
rect -960 319288 3299 319290
rect -960 319232 3238 319288
rect 3294 319232 3299 319288
rect -960 319230 3299 319232
rect -960 319140 480 319230
rect 3233 319227 3299 319230
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 2865 228034 2931 228037
rect -960 228032 2931 228034
rect -960 227976 2870 228032
rect 2926 227976 2931 228032
rect -960 227974 2931 227976
rect -960 227884 480 227974
rect 2865 227971 2931 227974
rect 580073 219058 580139 219061
rect 583520 219058 584960 219148
rect 580073 219056 584960 219058
rect 580073 219000 580078 219056
rect 580134 219000 584960 219056
rect 580073 218998 584960 219000
rect 580073 218995 580139 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580073 205730 580139 205733
rect 583520 205730 584960 205820
rect 580073 205728 584960 205730
rect 580073 205672 580078 205728
rect 580134 205672 584960 205728
rect 580073 205670 584960 205672
rect 580073 205667 580139 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 160093 195938 160159 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 158854 195936 160159 195938
rect 158854 195933 160098 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 158805 195928 160098 195933
rect 158805 195872 158810 195928
rect 158866 195880 160098 195928
rect 160154 195880 160159 195936
rect 158866 195878 160159 195880
rect 158866 195872 158914 195878
rect 160093 195875 160159 195878
rect 158805 195870 158914 195872
rect 158805 195867 158871 195870
rect 140773 195666 140839 195669
rect 143582 195666 144164 195674
rect 140773 195664 144164 195666
rect 140773 195608 140778 195664
rect 140834 195614 144164 195664
rect 140834 195608 143642 195614
rect 140773 195606 143642 195608
rect 140773 195603 140839 195606
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 579797 192538 579863 192541
rect 583520 192538 584960 192628
rect 579797 192536 584960 192538
rect 579797 192480 579802 192536
rect 579858 192480 584960 192536
rect 579797 192478 584960 192480
rect 579797 192475 579863 192478
rect 583520 192388 584960 192478
rect 140865 191858 140931 191861
rect 143582 191858 143980 191900
rect 140865 191856 143980 191858
rect 140865 191800 140870 191856
rect 140926 191840 143980 191856
rect 140926 191800 143642 191840
rect 140865 191798 143642 191800
rect 140865 191795 140931 191798
rect 140773 191586 140839 191589
rect 143582 191586 144164 191630
rect 140773 191584 144164 191586
rect 140773 191528 140778 191584
rect 140834 191570 144164 191584
rect 140834 191528 143642 191570
rect 140773 191526 143642 191528
rect 140773 191523 140839 191526
rect 140957 190906 141023 190909
rect 144134 190906 144194 191460
rect 144361 191042 144427 191045
rect 144494 191042 144500 191044
rect 144361 191040 144500 191042
rect 144361 190984 144366 191040
rect 144422 190984 144500 191040
rect 144361 190982 144500 190984
rect 144361 190979 144427 190982
rect 144494 190980 144500 190982
rect 144564 190980 144570 191044
rect 140957 190904 144194 190906
rect 140957 190848 140962 190904
rect 141018 190848 144194 190904
rect 140957 190846 144194 190848
rect 140957 190843 141023 190846
rect 145833 189000 145899 189005
rect -960 188866 480 188956
rect 145833 188944 145838 189000
rect 145894 188944 145899 189000
rect 145833 188939 145899 188944
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 145836 188594 145896 188939
rect 146150 188594 146156 188596
rect 145836 188534 146156 188594
rect 146150 188532 146156 188534
rect 146220 188532 146226 188596
rect 144494 188124 144500 188188
rect 144564 188186 144570 188188
rect 144913 188186 144979 188189
rect 144564 188184 144979 188186
rect 144564 188128 144918 188184
rect 144974 188128 144979 188184
rect 144564 188126 144979 188128
rect 144564 188124 144570 188126
rect 144913 188123 144979 188126
rect 140865 184378 140931 184381
rect 141182 184378 141188 184380
rect 140865 184376 141188 184378
rect 140865 184320 140870 184376
rect 140926 184320 141188 184376
rect 140865 184318 141188 184320
rect 140865 184315 140931 184318
rect 141182 184316 141188 184318
rect 141252 184316 141258 184380
rect 140773 184242 140839 184245
rect 140998 184242 141004 184244
rect 140773 184240 141004 184242
rect 140773 184184 140778 184240
rect 140834 184184 141004 184240
rect 140773 184182 141004 184184
rect 140773 184179 140839 184182
rect 140998 184180 141004 184182
rect 141068 184180 141074 184244
rect 140957 184106 141023 184109
rect 143022 184106 143028 184108
rect 140957 184104 143028 184106
rect 140957 184048 140962 184104
rect 141018 184048 143028 184104
rect 140957 184046 143028 184048
rect 140957 184043 141023 184046
rect 143022 184044 143028 184046
rect 143092 184044 143098 184108
rect 144913 181250 144979 181253
rect 148726 181250 148732 181252
rect 144913 181248 148732 181250
rect 144913 181192 144918 181248
rect 144974 181192 148732 181248
rect 144913 181190 148732 181192
rect 144913 181187 144979 181190
rect 148726 181188 148732 181190
rect 148796 181188 148802 181252
rect 144637 180980 144703 180981
rect 144637 180976 144684 180980
rect 144748 180978 144754 180980
rect 144637 180920 144642 180976
rect 144637 180916 144684 180920
rect 144748 180918 144794 180978
rect 144748 180916 144754 180918
rect 144637 180915 144703 180916
rect 157793 179482 157859 179485
rect 158529 179482 158595 179485
rect 157793 179480 158595 179482
rect 157793 179424 157798 179480
rect 157854 179424 158534 179480
rect 158590 179424 158595 179480
rect 157793 179422 158595 179424
rect 157793 179419 157859 179422
rect 158529 179419 158595 179422
rect 580073 179210 580139 179213
rect 583520 179210 584960 179300
rect 580073 179208 584960 179210
rect 580073 179152 580078 179208
rect 580134 179152 584960 179208
rect 580073 179150 584960 179152
rect 580073 179147 580139 179150
rect 583520 179060 584960 179150
rect 143022 178876 143028 178940
rect 143092 178938 143098 178940
rect 144085 178938 144151 178941
rect 143092 178936 144151 178938
rect 143092 178880 144090 178936
rect 144146 178880 144151 178936
rect 143092 178878 144151 178880
rect 143092 178876 143098 178878
rect 144085 178875 144151 178878
rect 141182 178740 141188 178804
rect 141252 178802 141258 178804
rect 143073 178802 143139 178805
rect 141252 178800 143139 178802
rect 141252 178744 143078 178800
rect 143134 178744 143139 178800
rect 141252 178742 143139 178744
rect 141252 178740 141258 178742
rect 143073 178739 143139 178742
rect 140998 178604 141004 178668
rect 141068 178666 141074 178668
rect 141601 178666 141667 178669
rect 141068 178664 141667 178666
rect 141068 178608 141606 178664
rect 141662 178608 141667 178664
rect 141068 178606 141667 178608
rect 141068 178604 141074 178606
rect 141601 178603 141667 178606
rect -960 175796 480 176036
rect 163497 175946 163563 175949
rect 165153 175946 165219 175949
rect 163497 175944 165219 175946
rect 163497 175888 163502 175944
rect 163558 175888 165158 175944
rect 165214 175888 165219 175944
rect 163497 175886 165219 175888
rect 163497 175883 163563 175886
rect 165153 175883 165219 175886
rect 163589 175810 163655 175813
rect 165061 175810 165127 175813
rect 163589 175808 165127 175810
rect 163589 175752 163594 175808
rect 163650 175752 165066 175808
rect 165122 175752 165127 175808
rect 163589 175750 165127 175752
rect 163589 175747 163655 175750
rect 165061 175747 165127 175750
rect 149329 175674 149395 175677
rect 158161 175674 158227 175677
rect 149329 175672 158227 175674
rect 149329 175616 149334 175672
rect 149390 175616 158166 175672
rect 158222 175616 158227 175672
rect 149329 175614 158227 175616
rect 149329 175611 149395 175614
rect 158161 175611 158227 175614
rect 148726 171804 148732 171868
rect 148796 171866 148802 171868
rect 155217 171866 155283 171869
rect 148796 171864 155283 171866
rect 148796 171808 155222 171864
rect 155278 171808 155283 171864
rect 148796 171806 155283 171808
rect 148796 171804 148802 171806
rect 155217 171803 155283 171806
rect 580073 165882 580139 165885
rect 583520 165882 584960 165972
rect 580073 165880 584960 165882
rect 580073 165824 580078 165880
rect 580134 165824 584960 165880
rect 580073 165822 584960 165824
rect 580073 165819 580139 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 4061 149834 4127 149837
rect -960 149832 4127 149834
rect -960 149776 4066 149832
rect 4122 149776 4127 149832
rect -960 149774 4127 149776
rect -960 149684 480 149774
rect 4061 149771 4127 149774
rect 146150 142836 146156 142900
rect 146220 142898 146226 142900
rect 171501 142898 171567 142901
rect 146220 142896 171567 142898
rect 146220 142840 171506 142896
rect 171562 142840 171567 142896
rect 146220 142838 171567 142840
rect 146220 142836 146226 142838
rect 171501 142835 171567 142838
rect 144678 142700 144684 142764
rect 144748 142762 144754 142764
rect 173065 142762 173131 142765
rect 144748 142760 173131 142762
rect 144748 142704 173070 142760
rect 173126 142704 173131 142760
rect 144748 142702 173131 142704
rect 144748 142700 144754 142702
rect 173065 142699 173131 142702
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 121269 138954 121335 138957
rect 120582 138952 121335 138954
rect 120582 138896 121274 138952
rect 121330 138896 121335 138952
rect 120582 138894 121335 138896
rect 120582 138380 120642 138894
rect 121269 138891 121335 138894
rect 180885 137594 180951 137597
rect 179860 137592 180951 137594
rect 179860 137536 180890 137592
rect 180946 137536 180951 137592
rect 179860 137534 180951 137536
rect 180885 137531 180951 137534
rect 117313 136914 117379 136917
rect 117313 136912 120060 136914
rect -960 136778 480 136868
rect 117313 136856 117318 136912
rect 117374 136856 120060 136912
rect 117313 136854 120060 136856
rect 117313 136851 117379 136854
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 179646 135557 179706 136068
rect 179597 135552 179706 135557
rect 179597 135496 179602 135552
rect 179658 135496 179706 135552
rect 179597 135494 179706 135496
rect 179597 135491 179663 135494
rect 117313 135418 117379 135421
rect 117313 135416 120060 135418
rect 117313 135360 117318 135416
rect 117374 135360 120060 135416
rect 117313 135358 120060 135360
rect 117313 135355 117379 135358
rect 182173 134602 182239 134605
rect 179860 134600 182239 134602
rect 179860 134544 182178 134600
rect 182234 134544 182239 134600
rect 179860 134542 182239 134544
rect 182173 134539 182239 134542
rect 117313 133922 117379 133925
rect 117313 133920 120060 133922
rect 117313 133864 117318 133920
rect 117374 133864 120060 133920
rect 117313 133862 120060 133864
rect 117313 133859 117379 133862
rect 181253 133106 181319 133109
rect 179860 133104 181319 133106
rect 179860 133048 181258 133104
rect 181314 133048 181319 133104
rect 179860 133046 181319 133048
rect 181253 133043 181319 133046
rect 117313 132426 117379 132429
rect 117313 132424 120060 132426
rect 117313 132368 117318 132424
rect 117374 132368 120060 132424
rect 117313 132366 120060 132368
rect 117313 132363 117379 132366
rect 179505 132018 179571 132021
rect 179462 132016 179571 132018
rect 179462 131960 179510 132016
rect 179566 131960 179571 132016
rect 179462 131955 179571 131960
rect 179462 131580 179522 131955
rect 117313 130930 117379 130933
rect 117313 130928 120060 130930
rect 117313 130872 117318 130928
rect 117374 130872 120060 130928
rect 117313 130870 120060 130872
rect 117313 130867 117379 130870
rect 182909 130114 182975 130117
rect 179860 130112 182975 130114
rect 179860 130056 182914 130112
rect 182970 130056 182975 130112
rect 179860 130054 182975 130056
rect 182909 130051 182975 130054
rect 117313 129434 117379 129437
rect 117313 129432 120060 129434
rect 117313 129376 117318 129432
rect 117374 129376 120060 129432
rect 117313 129374 120060 129376
rect 117313 129371 117379 129374
rect 182633 128618 182699 128621
rect 179860 128616 182699 128618
rect 179860 128560 182638 128616
rect 182694 128560 182699 128616
rect 179860 128558 182699 128560
rect 182633 128555 182699 128558
rect 117313 127938 117379 127941
rect 117313 127936 120060 127938
rect 117313 127880 117318 127936
rect 117374 127880 120060 127936
rect 117313 127878 120060 127880
rect 117313 127875 117379 127878
rect 182541 127122 182607 127125
rect 179860 127120 182607 127122
rect 179860 127064 182546 127120
rect 182602 127064 182607 127120
rect 179860 127062 182607 127064
rect 182541 127059 182607 127062
rect 117313 126442 117379 126445
rect 117313 126440 120060 126442
rect 117313 126384 117318 126440
rect 117374 126384 120060 126440
rect 117313 126382 120060 126384
rect 117313 126379 117379 126382
rect 179413 126170 179479 126173
rect 179413 126168 179522 126170
rect 179413 126112 179418 126168
rect 179474 126112 179522 126168
rect 179413 126107 179522 126112
rect 179462 125596 179522 126107
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 117313 124946 117379 124949
rect 117313 124944 120060 124946
rect 117313 124888 117318 124944
rect 117374 124888 120060 124944
rect 117313 124886 120060 124888
rect 117313 124883 117379 124886
rect 180793 124130 180859 124133
rect 179860 124128 180859 124130
rect 179860 124072 180798 124128
rect 180854 124072 180859 124128
rect 179860 124070 180859 124072
rect 180793 124067 180859 124070
rect -960 123572 480 123812
rect 117313 123450 117379 123453
rect 117313 123448 120060 123450
rect 117313 123392 117318 123448
rect 117374 123392 120060 123448
rect 117313 123390 120060 123392
rect 117313 123387 117379 123390
rect 182265 122634 182331 122637
rect 179860 122632 182331 122634
rect 179860 122576 182270 122632
rect 182326 122576 182331 122632
rect 179860 122574 182331 122576
rect 182265 122571 182331 122574
rect 117313 121954 117379 121957
rect 117313 121952 120060 121954
rect 117313 121896 117318 121952
rect 117374 121896 120060 121952
rect 117313 121894 120060 121896
rect 117313 121891 117379 121894
rect 182725 121138 182791 121141
rect 179860 121136 182791 121138
rect 179860 121080 182730 121136
rect 182786 121080 182791 121136
rect 179860 121078 182791 121080
rect 182725 121075 182791 121078
rect 117313 120458 117379 120461
rect 117313 120456 120060 120458
rect 117313 120400 117318 120456
rect 117374 120400 120060 120456
rect 117313 120398 120060 120400
rect 117313 120395 117379 120398
rect 182449 119642 182515 119645
rect 179860 119640 182515 119642
rect 179860 119584 182454 119640
rect 182510 119584 182515 119640
rect 179860 119582 182515 119584
rect 182449 119579 182515 119582
rect 117313 118962 117379 118965
rect 117313 118960 120060 118962
rect 117313 118904 117318 118960
rect 117374 118904 120060 118960
rect 117313 118902 120060 118904
rect 117313 118899 117379 118902
rect 182357 118146 182423 118149
rect 179860 118144 182423 118146
rect 179860 118088 182362 118144
rect 182418 118088 182423 118144
rect 179860 118086 182423 118088
rect 182357 118083 182423 118086
rect 117313 117466 117379 117469
rect 117313 117464 120060 117466
rect 117313 117408 117318 117464
rect 117374 117408 120060 117464
rect 117313 117406 120060 117408
rect 117313 117403 117379 117406
rect 180977 116650 181043 116653
rect 179860 116648 181043 116650
rect 179860 116592 180982 116648
rect 181038 116592 181043 116648
rect 179860 116590 181043 116592
rect 180977 116587 181043 116590
rect 117313 115970 117379 115973
rect 117313 115968 120060 115970
rect 117313 115912 117318 115968
rect 117374 115912 120060 115968
rect 117313 115910 120060 115912
rect 117313 115907 117379 115910
rect 181161 115154 181227 115157
rect 179860 115152 181227 115154
rect 179860 115096 181166 115152
rect 181222 115096 181227 115152
rect 179860 115094 181227 115096
rect 181161 115091 181227 115094
rect 117313 114474 117379 114477
rect 117313 114472 120060 114474
rect 117313 114416 117318 114472
rect 117374 114416 120060 114472
rect 117313 114414 120060 114416
rect 117313 114411 117379 114414
rect 182173 113658 182239 113661
rect 179860 113656 182239 113658
rect 179860 113600 182178 113656
rect 182234 113600 182239 113656
rect 179860 113598 182239 113600
rect 182173 113595 182239 113598
rect 117313 112978 117379 112981
rect 117313 112976 120060 112978
rect 117313 112920 117318 112976
rect 117374 112920 120060 112976
rect 117313 112918 120060 112920
rect 117313 112915 117379 112918
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 181069 112162 181135 112165
rect 179860 112160 181135 112162
rect 179860 112104 181074 112160
rect 181130 112104 181135 112160
rect 179860 112102 181135 112104
rect 181069 112099 181135 112102
rect 117313 111482 117379 111485
rect 117313 111480 120060 111482
rect 117313 111424 117318 111480
rect 117374 111424 120060 111480
rect 117313 111422 120060 111424
rect 117313 111419 117379 111422
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect 183277 110666 183343 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect 179860 110664 183343 110666
rect 179860 110608 183282 110664
rect 183338 110608 183343 110664
rect 179860 110606 183343 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 183277 110603 183343 110606
rect 117313 109986 117379 109989
rect 117313 109984 120060 109986
rect 117313 109928 117318 109984
rect 117374 109928 120060 109984
rect 117313 109926 120060 109928
rect 117313 109923 117379 109926
rect 183461 109170 183527 109173
rect 179860 109168 183527 109170
rect 179860 109112 183466 109168
rect 183522 109112 183527 109168
rect 179860 109110 183527 109112
rect 183461 109107 183527 109110
rect 118049 108490 118115 108493
rect 118049 108488 120060 108490
rect 118049 108432 118054 108488
rect 118110 108432 120060 108488
rect 118049 108430 120060 108432
rect 118049 108427 118115 108430
rect 183369 107674 183435 107677
rect 179860 107672 183435 107674
rect 179860 107616 183374 107672
rect 183430 107616 183435 107672
rect 179860 107614 183435 107616
rect 183369 107611 183435 107614
rect 117865 106994 117931 106997
rect 117865 106992 120060 106994
rect 117865 106936 117870 106992
rect 117926 106936 120060 106992
rect 117865 106934 120060 106936
rect 117865 106931 117931 106934
rect 183461 106178 183527 106181
rect 179860 106176 183527 106178
rect 179860 106120 183466 106176
rect 183522 106120 183527 106176
rect 179860 106118 183527 106120
rect 183461 106115 183527 106118
rect 120625 106042 120691 106045
rect 120582 106040 120691 106042
rect 120582 105984 120630 106040
rect 120686 105984 120691 106040
rect 120582 105979 120691 105984
rect 120582 105468 120642 105979
rect 183461 104682 183527 104685
rect 179860 104680 183527 104682
rect 179860 104624 183466 104680
rect 183522 104624 183527 104680
rect 179860 104622 183527 104624
rect 183461 104619 183527 104622
rect 118141 104002 118207 104005
rect 118141 104000 120060 104002
rect 118141 103944 118146 104000
rect 118202 103944 120060 104000
rect 118141 103942 120060 103944
rect 118141 103939 118207 103942
rect 183461 103186 183527 103189
rect 179860 103184 183527 103186
rect 179860 103128 183466 103184
rect 183522 103128 183527 103184
rect 179860 103126 183527 103128
rect 183461 103123 183527 103126
rect 119245 102506 119311 102509
rect 119245 102504 120060 102506
rect 119245 102448 119250 102504
rect 119306 102448 120060 102504
rect 119245 102446 120060 102448
rect 119245 102443 119311 102446
rect 183461 101690 183527 101693
rect 179860 101688 183527 101690
rect 179860 101632 183466 101688
rect 183522 101632 183527 101688
rect 179860 101630 183527 101632
rect 183461 101627 183527 101630
rect 118785 101010 118851 101013
rect 118785 101008 120060 101010
rect 118785 100952 118790 101008
rect 118846 100952 120060 101008
rect 118785 100950 120060 100952
rect 118785 100947 118851 100950
rect 183461 100194 183527 100197
rect 179860 100192 183527 100194
rect 179860 100136 183466 100192
rect 183522 100136 183527 100192
rect 179860 100134 183527 100136
rect 183461 100131 183527 100134
rect 119153 99514 119219 99517
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 119153 99512 120060 99514
rect 119153 99456 119158 99512
rect 119214 99456 120060 99512
rect 119153 99454 120060 99456
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 119153 99451 119219 99454
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect 183461 98698 183527 98701
rect 179860 98696 183527 98698
rect 179860 98640 183466 98696
rect 183522 98640 183527 98696
rect 179860 98638 183527 98640
rect 183461 98635 183527 98638
rect 118969 98018 119035 98021
rect 118969 98016 120060 98018
rect 118969 97960 118974 98016
rect 119030 97960 120060 98016
rect 118969 97958 120060 97960
rect 118969 97955 119035 97958
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 183461 97202 183527 97205
rect 179860 97200 183527 97202
rect 179860 97144 183466 97200
rect 183522 97144 183527 97200
rect 179860 97142 183527 97144
rect 183461 97139 183527 97142
rect 119061 96522 119127 96525
rect 119061 96520 120060 96522
rect 119061 96464 119066 96520
rect 119122 96464 120060 96520
rect 119061 96462 120060 96464
rect 119061 96459 119127 96462
rect 183185 95706 183251 95709
rect 179860 95704 183251 95706
rect 179860 95648 183190 95704
rect 183246 95648 183251 95704
rect 179860 95646 183251 95648
rect 183185 95643 183251 95646
rect 118233 95026 118299 95029
rect 118233 95024 120060 95026
rect 118233 94968 118238 95024
rect 118294 94968 120060 95024
rect 118233 94966 120060 94968
rect 118233 94963 118299 94966
rect 183277 94210 183343 94213
rect 179860 94208 183343 94210
rect 179860 94152 183282 94208
rect 183338 94152 183343 94208
rect 179860 94150 183343 94152
rect 183277 94147 183343 94150
rect 118325 93530 118391 93533
rect 118325 93528 120060 93530
rect 118325 93472 118330 93528
rect 118386 93472 120060 93528
rect 118325 93470 120060 93472
rect 118325 93467 118391 93470
rect 183277 92714 183343 92717
rect 179860 92712 183343 92714
rect 179860 92656 183282 92712
rect 183338 92656 183343 92712
rect 179860 92654 183343 92656
rect 183277 92651 183343 92654
rect 118417 92034 118483 92037
rect 118417 92032 120060 92034
rect 118417 91976 118422 92032
rect 118478 91976 120060 92032
rect 118417 91974 120060 91976
rect 118417 91971 118483 91974
rect 183461 91218 183527 91221
rect 179860 91216 183527 91218
rect 179860 91160 183466 91216
rect 183522 91160 183527 91216
rect 179860 91158 183527 91160
rect 183461 91155 183527 91158
rect 118509 90538 118575 90541
rect 118509 90536 120060 90538
rect 118509 90480 118514 90536
rect 118570 90480 120060 90536
rect 118509 90478 120060 90480
rect 118509 90475 118575 90478
rect 183461 89722 183527 89725
rect 179860 89720 183527 89722
rect 179860 89664 183466 89720
rect 183522 89664 183527 89720
rect 179860 89662 183527 89664
rect 183461 89659 183527 89662
rect 118693 89042 118759 89045
rect 118693 89040 120060 89042
rect 118693 88984 118698 89040
rect 118754 88984 120060 89040
rect 118693 88982 120060 88984
rect 118693 88979 118759 88982
rect 183461 88226 183527 88229
rect 179860 88224 183527 88226
rect 179860 88168 183466 88224
rect 183522 88168 183527 88224
rect 179860 88166 183527 88168
rect 183461 88163 183527 88166
rect 118877 87546 118943 87549
rect 118877 87544 120060 87546
rect 118877 87488 118882 87544
rect 118938 87488 120060 87544
rect 118877 87486 120060 87488
rect 118877 87483 118943 87486
rect 182817 86730 182883 86733
rect 179860 86728 182883 86730
rect 179860 86672 182822 86728
rect 182878 86672 182883 86728
rect 179860 86670 182883 86672
rect 182817 86667 182883 86670
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 118601 86050 118667 86053
rect 118601 86048 120060 86050
rect 118601 85992 118606 86048
rect 118662 85992 120060 86048
rect 583520 86036 584960 86126
rect 118601 85990 120060 85992
rect 118601 85987 118667 85990
rect 183461 85234 183527 85237
rect 179860 85232 183527 85234
rect 179860 85176 183466 85232
rect 183522 85176 183527 85232
rect 179860 85174 183527 85176
rect 183461 85171 183527 85174
rect -960 84690 480 84780
rect 3969 84690 4035 84693
rect -960 84688 4035 84690
rect -960 84632 3974 84688
rect 4030 84632 4035 84688
rect -960 84630 4035 84632
rect -960 84540 480 84630
rect 3969 84627 4035 84630
rect 120582 84285 120642 84524
rect 120582 84280 120691 84285
rect 120582 84224 120630 84280
rect 120686 84224 120691 84280
rect 120582 84222 120691 84224
rect 120625 84219 120691 84222
rect 182817 83738 182883 83741
rect 179860 83736 182883 83738
rect 179860 83680 182822 83736
rect 182878 83680 182883 83736
rect 179860 83678 182883 83680
rect 182817 83675 182883 83678
rect 118509 83058 118575 83061
rect 118509 83056 120060 83058
rect 118509 83000 118514 83056
rect 118570 83000 120060 83056
rect 118509 82998 120060 83000
rect 118509 82995 118575 82998
rect 183461 82242 183527 82245
rect 179860 82240 183527 82242
rect 179860 82184 183466 82240
rect 183522 82184 183527 82240
rect 179860 82182 183527 82184
rect 183461 82179 183527 82182
rect 118417 81562 118483 81565
rect 118417 81560 120060 81562
rect 118417 81504 118422 81560
rect 118478 81504 120060 81560
rect 118417 81502 120060 81504
rect 118417 81499 118483 81502
rect 120625 81426 120691 81429
rect 580257 81426 580323 81429
rect 120625 81424 580323 81426
rect 120625 81368 120630 81424
rect 120686 81368 580262 81424
rect 580318 81368 580323 81424
rect 120625 81366 580323 81368
rect 120625 81363 120691 81366
rect 580257 81363 580323 81366
rect 3509 81290 3575 81293
rect 173382 81290 173388 81292
rect 3509 81288 173388 81290
rect 3509 81232 3514 81288
rect 3570 81232 173388 81288
rect 3509 81230 173388 81232
rect 3509 81227 3575 81230
rect 173382 81228 173388 81230
rect 173452 81228 173458 81292
rect 180057 81290 180123 81293
rect 173528 81288 180123 81290
rect 173528 81232 180062 81288
rect 180118 81232 180123 81288
rect 173528 81230 180123 81232
rect 171174 81092 171180 81156
rect 171244 81154 171250 81156
rect 173528 81154 173588 81230
rect 180057 81227 180123 81230
rect 396809 81154 396875 81157
rect 171244 81094 173588 81154
rect 173666 81152 396875 81154
rect 173666 81096 396814 81152
rect 396870 81096 396875 81152
rect 173666 81094 396875 81096
rect 171244 81092 171250 81094
rect 171910 80956 171916 81020
rect 171980 81018 171986 81020
rect 173666 81018 173726 81094
rect 396809 81091 396875 81094
rect 171980 80958 173726 81018
rect 178401 81018 178467 81021
rect 396993 81018 397059 81021
rect 178401 81016 397059 81018
rect 178401 80960 178406 81016
rect 178462 80960 396998 81016
rect 397054 80960 397059 81016
rect 178401 80958 397059 80960
rect 171980 80956 171986 80958
rect 178401 80955 178467 80958
rect 396993 80955 397059 80958
rect 178309 80882 178375 80885
rect 504357 80882 504423 80885
rect 178309 80880 504423 80882
rect 178309 80824 178314 80880
rect 178370 80824 504362 80880
rect 504418 80824 504423 80880
rect 178309 80822 504423 80824
rect 178309 80819 178375 80822
rect 504357 80819 504423 80822
rect 172094 80684 172100 80748
rect 172164 80746 172170 80748
rect 580901 80746 580967 80749
rect 172164 80744 580967 80746
rect 172164 80688 580906 80744
rect 580962 80688 580967 80744
rect 172164 80686 580967 80688
rect 172164 80684 172170 80686
rect 580901 80683 580967 80686
rect 3877 80610 3943 80613
rect 173014 80610 173020 80612
rect 3877 80608 173020 80610
rect 3877 80552 3882 80608
rect 3938 80552 173020 80608
rect 3877 80550 173020 80552
rect 3877 80547 3943 80550
rect 173014 80548 173020 80550
rect 173084 80548 173090 80612
rect 3141 80474 3207 80477
rect 172830 80474 172836 80476
rect 3141 80472 172836 80474
rect 3141 80416 3146 80472
rect 3202 80416 172836 80472
rect 3141 80414 172836 80416
rect 3141 80411 3207 80414
rect 172830 80412 172836 80414
rect 172900 80412 172906 80476
rect 171358 80338 171364 80340
rect 163224 80278 171364 80338
rect 158662 80140 158668 80204
rect 158732 80202 158738 80204
rect 158732 80142 159006 80202
rect 158732 80140 158738 80142
rect 130326 80066 130332 80068
rect 130058 80006 130332 80066
rect 126375 79964 126441 79967
rect 127111 79964 127177 79967
rect 126375 79962 126484 79964
rect 125731 79932 125797 79933
rect 125726 79868 125732 79932
rect 125796 79930 125802 79932
rect 125796 79870 125888 79930
rect 126099 79928 126165 79933
rect 126099 79872 126104 79928
rect 126160 79872 126165 79928
rect 126375 79906 126380 79962
rect 126436 79906 126484 79962
rect 127068 79962 127177 79964
rect 127068 79932 127116 79962
rect 126375 79901 126484 79906
rect 125796 79868 125802 79870
rect 125731 79867 125797 79868
rect 126099 79867 126165 79872
rect 123017 79794 123083 79797
rect 126102 79794 126162 79867
rect 123017 79792 126162 79794
rect 123017 79736 123022 79792
rect 123078 79736 126162 79792
rect 123017 79734 126162 79736
rect 123017 79731 123083 79734
rect 126145 79658 126211 79661
rect 126424 79658 126484 79901
rect 127014 79868 127020 79932
rect 127084 79906 127116 79932
rect 127172 79906 127177 79962
rect 127847 79964 127913 79967
rect 127847 79962 127956 79964
rect 127084 79901 127177 79906
rect 127295 79930 127361 79933
rect 127295 79928 127588 79930
rect 127084 79870 127128 79901
rect 127295 79872 127300 79928
rect 127356 79872 127588 79928
rect 127847 79906 127852 79962
rect 127908 79906 127956 79962
rect 127847 79901 127956 79906
rect 128123 79962 128189 79967
rect 128123 79906 128128 79962
rect 128184 79906 128189 79962
rect 128123 79901 128189 79906
rect 128491 79962 128557 79967
rect 128491 79906 128496 79962
rect 128552 79906 128557 79962
rect 128675 79962 128741 79967
rect 128675 79932 128680 79962
rect 128736 79932 128741 79962
rect 128859 79962 128925 79967
rect 128491 79901 128557 79906
rect 127295 79870 127588 79872
rect 127084 79868 127090 79870
rect 127295 79867 127361 79870
rect 127198 79732 127204 79796
rect 127268 79794 127274 79796
rect 127528 79794 127588 79870
rect 127268 79734 127588 79794
rect 127709 79794 127775 79797
rect 127896 79794 127956 79901
rect 127709 79792 127956 79794
rect 127709 79736 127714 79792
rect 127770 79736 127956 79792
rect 127709 79734 127956 79736
rect 127268 79732 127274 79734
rect 127709 79731 127775 79734
rect 126145 79656 126484 79658
rect 126145 79600 126150 79656
rect 126206 79600 126484 79656
rect 126145 79598 126484 79600
rect 127525 79658 127591 79661
rect 128126 79658 128186 79901
rect 127525 79656 128186 79658
rect 127525 79600 127530 79656
rect 127586 79600 128186 79656
rect 127525 79598 128186 79600
rect 128494 79658 128554 79901
rect 128670 79868 128676 79932
rect 128740 79930 128746 79932
rect 128740 79870 128798 79930
rect 128859 79906 128864 79962
rect 128920 79906 128925 79962
rect 130058 79933 130118 80006
rect 130326 80004 130332 80006
rect 130396 80004 130402 80068
rect 144678 80004 144684 80068
rect 144748 80066 144754 80068
rect 144748 80004 144792 80066
rect 151486 80004 151492 80068
rect 151556 80004 151562 80068
rect 131251 79962 131317 79967
rect 128859 79901 128925 79906
rect 129227 79928 129293 79933
rect 128740 79868 128746 79870
rect 128862 79796 128922 79901
rect 129227 79872 129232 79928
rect 129288 79872 129293 79928
rect 129227 79867 129293 79872
rect 130055 79928 130121 79933
rect 130055 79872 130060 79928
rect 130116 79872 130121 79928
rect 130055 79867 130121 79872
rect 130331 79930 130397 79933
rect 131251 79932 131256 79962
rect 131312 79932 131317 79962
rect 131435 79962 131501 79967
rect 130510 79930 130516 79932
rect 130331 79928 130516 79930
rect 130331 79872 130336 79928
rect 130392 79872 130516 79928
rect 130331 79870 130516 79872
rect 130331 79867 130397 79870
rect 130510 79868 130516 79870
rect 130580 79868 130586 79932
rect 131246 79868 131252 79932
rect 131316 79930 131322 79932
rect 131316 79870 131374 79930
rect 131435 79906 131440 79962
rect 131496 79906 131501 79962
rect 131619 79962 131685 79967
rect 131619 79932 131624 79962
rect 131680 79932 131685 79962
rect 131895 79964 131961 79967
rect 131895 79962 132234 79964
rect 131435 79901 131501 79906
rect 131316 79868 131322 79870
rect 128854 79732 128860 79796
rect 128924 79732 128930 79796
rect 129230 79661 129290 79867
rect 131438 79797 131498 79901
rect 131614 79868 131620 79932
rect 131684 79930 131690 79932
rect 131684 79870 131742 79930
rect 131895 79906 131900 79962
rect 131956 79906 132234 79962
rect 131895 79904 132234 79906
rect 131895 79901 131961 79904
rect 131684 79868 131690 79870
rect 131389 79792 131498 79797
rect 131389 79736 131394 79792
rect 131450 79736 131498 79792
rect 131389 79734 131498 79736
rect 131389 79731 131455 79734
rect 129038 79658 129044 79660
rect 128494 79598 129044 79658
rect 126145 79595 126211 79598
rect 127525 79595 127591 79598
rect 129038 79596 129044 79598
rect 129108 79596 129114 79660
rect 129181 79656 129290 79661
rect 129181 79600 129186 79656
rect 129242 79600 129290 79656
rect 129181 79598 129290 79600
rect 131849 79658 131915 79661
rect 132174 79658 132234 79904
rect 132355 79962 132421 79967
rect 132355 79906 132360 79962
rect 132416 79906 132421 79962
rect 132355 79901 132421 79906
rect 132631 79962 132697 79967
rect 132631 79906 132636 79962
rect 132692 79930 132697 79962
rect 134195 79962 134261 79967
rect 133270 79930 133276 79932
rect 132692 79906 133276 79930
rect 132631 79901 133276 79906
rect 132358 79797 132418 79901
rect 132634 79870 133276 79901
rect 133270 79868 133276 79870
rect 133340 79868 133346 79932
rect 133827 79930 133893 79933
rect 134195 79932 134200 79962
rect 134256 79932 134261 79962
rect 134379 79962 134445 79967
rect 133646 79928 133893 79930
rect 133459 79894 133525 79899
rect 133459 79838 133464 79894
rect 133520 79838 133525 79894
rect 133459 79833 133525 79838
rect 133646 79872 133832 79928
rect 133888 79872 133893 79928
rect 133646 79870 133893 79872
rect 132309 79792 132418 79797
rect 132309 79736 132314 79792
rect 132370 79736 132418 79792
rect 132309 79734 132418 79736
rect 132309 79731 132375 79734
rect 131849 79656 132234 79658
rect 131849 79600 131854 79656
rect 131910 79600 132234 79656
rect 131849 79598 132234 79600
rect 132493 79658 132559 79661
rect 133462 79658 133522 79833
rect 132493 79656 133522 79658
rect 132493 79600 132498 79656
rect 132554 79600 133522 79656
rect 132493 79598 133522 79600
rect 133646 79658 133706 79870
rect 133827 79867 133893 79870
rect 134190 79868 134196 79932
rect 134260 79930 134266 79932
rect 134260 79870 134318 79930
rect 134379 79906 134384 79962
rect 134440 79906 134445 79962
rect 136035 79962 136101 79967
rect 134839 79930 134905 79933
rect 135391 79930 135457 79933
rect 135759 79930 135825 79933
rect 134379 79901 134445 79906
rect 134566 79928 134905 79930
rect 134260 79868 134266 79870
rect 134382 79797 134442 79901
rect 134011 79796 134077 79797
rect 134006 79794 134012 79796
rect 133920 79734 134012 79794
rect 134006 79732 134012 79734
rect 134076 79732 134082 79796
rect 134333 79792 134442 79797
rect 134333 79736 134338 79792
rect 134394 79736 134442 79792
rect 134333 79734 134442 79736
rect 134566 79872 134844 79928
rect 134900 79872 134905 79928
rect 134566 79870 134905 79872
rect 134566 79794 134626 79870
rect 134839 79867 134905 79870
rect 135256 79928 135457 79930
rect 135256 79872 135396 79928
rect 135452 79872 135457 79928
rect 135256 79870 135457 79872
rect 134793 79794 134859 79797
rect 134566 79792 134859 79794
rect 134566 79736 134798 79792
rect 134854 79736 134859 79792
rect 134566 79734 134859 79736
rect 135256 79796 135316 79870
rect 135391 79867 135457 79870
rect 135578 79928 135825 79930
rect 135578 79872 135764 79928
rect 135820 79872 135825 79928
rect 136035 79906 136040 79962
rect 136096 79906 136101 79962
rect 136035 79901 136101 79906
rect 137139 79962 137205 79967
rect 137139 79906 137144 79962
rect 137200 79906 137205 79962
rect 137139 79901 137205 79906
rect 137323 79962 137389 79967
rect 137323 79906 137328 79962
rect 137384 79906 137389 79962
rect 138427 79964 138493 79967
rect 139991 79964 140057 79967
rect 141095 79964 141161 79967
rect 142015 79964 142081 79967
rect 138427 79962 138550 79964
rect 138427 79932 138432 79962
rect 138488 79932 138550 79962
rect 139991 79962 140192 79964
rect 137323 79901 137389 79906
rect 135578 79870 135825 79872
rect 135256 79734 135300 79796
rect 134011 79731 134077 79732
rect 134333 79731 134399 79734
rect 134793 79731 134859 79734
rect 135294 79732 135300 79734
rect 135364 79732 135370 79796
rect 135578 79794 135638 79870
rect 135759 79867 135825 79870
rect 135713 79794 135779 79797
rect 135578 79792 135779 79794
rect 135578 79736 135718 79792
rect 135774 79736 135779 79792
rect 135578 79734 135779 79736
rect 135713 79731 135779 79734
rect 136038 79661 136098 79901
rect 137142 79797 137202 79901
rect 137142 79792 137251 79797
rect 137142 79736 137190 79792
rect 137246 79736 137251 79792
rect 137142 79734 137251 79736
rect 137326 79794 137386 79901
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 137756 79870 138076 79930
rect 137756 79868 137762 79870
rect 138016 79797 138076 79870
rect 138422 79868 138428 79932
rect 138492 79904 138550 79932
rect 138979 79930 139045 79933
rect 139531 79930 139597 79933
rect 138614 79928 139045 79930
rect 138492 79868 138498 79904
rect 138614 79872 138984 79928
rect 139040 79872 139045 79928
rect 138614 79870 139045 79872
rect 137553 79794 137619 79797
rect 137326 79792 137619 79794
rect 137326 79736 137558 79792
rect 137614 79736 137619 79792
rect 137326 79734 137619 79736
rect 137185 79731 137251 79734
rect 137553 79731 137619 79734
rect 137967 79792 138076 79797
rect 138614 79796 138674 79870
rect 138979 79867 139045 79870
rect 139396 79928 139597 79930
rect 139396 79872 139536 79928
rect 139592 79872 139597 79928
rect 139991 79906 139996 79962
rect 140052 79906 140192 79962
rect 141095 79962 141204 79964
rect 139991 79904 140192 79906
rect 139991 79901 140057 79904
rect 139396 79870 139597 79872
rect 137967 79736 137972 79792
rect 138028 79736 138076 79792
rect 137967 79734 138076 79736
rect 137967 79731 138033 79734
rect 138606 79732 138612 79796
rect 138676 79732 138682 79796
rect 138974 79732 138980 79796
rect 139044 79794 139050 79796
rect 139163 79794 139229 79797
rect 139044 79792 139229 79794
rect 139044 79736 139168 79792
rect 139224 79736 139229 79792
rect 139044 79734 139229 79736
rect 139044 79732 139050 79734
rect 139163 79731 139229 79734
rect 139396 79661 139456 79870
rect 139531 79867 139597 79870
rect 139577 79794 139643 79797
rect 139945 79794 140011 79797
rect 139577 79792 140011 79794
rect 139577 79736 139582 79792
rect 139638 79736 139950 79792
rect 140006 79736 140011 79792
rect 139577 79734 140011 79736
rect 139577 79731 139643 79734
rect 139945 79731 140011 79734
rect 133781 79658 133847 79661
rect 133646 79656 133847 79658
rect 133646 79600 133786 79656
rect 133842 79600 133847 79656
rect 133646 79598 133847 79600
rect 129181 79595 129247 79598
rect 131849 79595 131915 79598
rect 132493 79595 132559 79598
rect 133781 79595 133847 79598
rect 134057 79658 134123 79661
rect 134190 79658 134196 79660
rect 134057 79656 134196 79658
rect 134057 79600 134062 79656
rect 134118 79600 134196 79656
rect 134057 79598 134196 79600
rect 134057 79595 134123 79598
rect 134190 79596 134196 79598
rect 134260 79596 134266 79660
rect 136038 79656 136147 79661
rect 136038 79600 136086 79656
rect 136142 79600 136147 79656
rect 136038 79598 136147 79600
rect 136081 79595 136147 79598
rect 139393 79656 139459 79661
rect 139393 79600 139398 79656
rect 139454 79600 139459 79656
rect 139393 79595 139459 79600
rect 139945 79658 140011 79661
rect 140132 79658 140192 79904
rect 140446 79868 140452 79932
rect 140516 79930 140522 79932
rect 140635 79930 140701 79933
rect 140516 79928 140701 79930
rect 140516 79872 140640 79928
rect 140696 79872 140701 79928
rect 141095 79906 141100 79962
rect 141156 79906 141204 79962
rect 141095 79901 141204 79906
rect 140516 79870 140701 79872
rect 140516 79868 140522 79870
rect 140635 79867 140701 79870
rect 141144 79794 141204 79901
rect 141972 79962 142081 79964
rect 141972 79906 142020 79962
rect 142076 79930 142081 79962
rect 142751 79964 142817 79967
rect 143303 79964 143369 79967
rect 142751 79962 142860 79964
rect 142470 79930 142476 79932
rect 142076 79906 142476 79930
rect 141972 79870 142476 79906
rect 142470 79868 142476 79870
rect 142540 79868 142546 79932
rect 142751 79906 142756 79962
rect 142812 79932 142860 79962
rect 143260 79962 143369 79964
rect 142812 79906 142844 79932
rect 142751 79901 142844 79906
rect 142800 79870 142844 79901
rect 142838 79868 142844 79870
rect 142908 79868 142914 79932
rect 143260 79906 143308 79962
rect 143364 79906 143369 79962
rect 143947 79962 144013 79967
rect 143487 79930 143553 79933
rect 143260 79901 143369 79906
rect 143444 79928 143553 79930
rect 142521 79794 142587 79797
rect 141144 79792 142587 79794
rect 141144 79736 142526 79792
rect 142582 79736 142587 79792
rect 141144 79734 142587 79736
rect 142521 79731 142587 79734
rect 142843 79792 142909 79797
rect 142843 79736 142848 79792
rect 142904 79736 142909 79792
rect 142843 79731 142909 79736
rect 143022 79732 143028 79796
rect 143092 79794 143098 79796
rect 143260 79794 143320 79901
rect 143092 79734 143320 79794
rect 143444 79872 143492 79928
rect 143548 79872 143553 79928
rect 143444 79867 143553 79872
rect 143758 79868 143764 79932
rect 143828 79930 143834 79932
rect 143947 79930 143952 79962
rect 143828 79906 143952 79930
rect 144008 79906 144013 79962
rect 143828 79901 144013 79906
rect 144315 79928 144381 79933
rect 143828 79870 144010 79901
rect 144315 79872 144320 79928
rect 144376 79872 144381 79928
rect 143828 79868 143834 79870
rect 144315 79867 144381 79872
rect 144591 79930 144657 79933
rect 144732 79930 144792 80004
rect 144591 79928 144792 79930
rect 144591 79872 144596 79928
rect 144652 79872 144792 79928
rect 144867 79962 144933 79967
rect 147351 79964 147417 79967
rect 144867 79906 144872 79962
rect 144928 79906 144933 79962
rect 147308 79962 147417 79964
rect 145511 79930 145577 79933
rect 145971 79932 146037 79933
rect 145966 79930 145972 79932
rect 144867 79901 144933 79906
rect 145238 79928 145577 79930
rect 144591 79870 144792 79872
rect 144591 79867 144657 79870
rect 143444 79794 143504 79867
rect 144126 79794 144132 79796
rect 143444 79734 144132 79794
rect 143092 79732 143098 79734
rect 144126 79732 144132 79734
rect 144196 79732 144202 79796
rect 142846 79661 142906 79731
rect 139945 79656 140192 79658
rect 139945 79600 139950 79656
rect 140006 79600 140192 79656
rect 139945 79598 140192 79600
rect 139945 79595 140011 79598
rect 140998 79596 141004 79660
rect 141068 79658 141074 79660
rect 142061 79658 142127 79661
rect 141068 79656 142127 79658
rect 141068 79600 142066 79656
rect 142122 79600 142127 79656
rect 141068 79598 142127 79600
rect 142846 79656 142955 79661
rect 143257 79660 143323 79661
rect 143206 79658 143212 79660
rect 142846 79600 142894 79656
rect 142950 79600 142955 79656
rect 142846 79598 142955 79600
rect 143166 79598 143212 79658
rect 143276 79656 143323 79660
rect 143318 79600 143323 79656
rect 141068 79596 141074 79598
rect 142061 79595 142127 79598
rect 142889 79595 142955 79598
rect 143206 79596 143212 79598
rect 143276 79596 143323 79600
rect 143257 79595 143323 79596
rect 143717 79658 143783 79661
rect 144318 79658 144378 79867
rect 144494 79732 144500 79796
rect 144564 79794 144570 79796
rect 144870 79794 144930 79901
rect 145051 79894 145117 79899
rect 145051 79838 145056 79894
rect 145112 79838 145117 79894
rect 145051 79833 145117 79838
rect 145238 79872 145516 79928
rect 145572 79872 145577 79928
rect 145238 79870 145577 79872
rect 145880 79870 145972 79930
rect 144564 79734 144930 79794
rect 144564 79732 144570 79734
rect 143717 79656 144378 79658
rect 143717 79600 143722 79656
rect 143778 79600 144378 79656
rect 143717 79598 144378 79600
rect 145054 79661 145114 79833
rect 145054 79656 145163 79661
rect 145054 79600 145102 79656
rect 145158 79600 145163 79656
rect 145054 79598 145163 79600
rect 145238 79658 145298 79870
rect 145511 79867 145577 79870
rect 145966 79868 145972 79870
rect 146036 79868 146042 79932
rect 146155 79930 146221 79933
rect 146112 79928 146221 79930
rect 146112 79872 146160 79928
rect 146216 79872 146221 79928
rect 145971 79867 146037 79868
rect 146112 79867 146221 79872
rect 146339 79928 146405 79933
rect 147308 79932 147356 79962
rect 146339 79872 146344 79928
rect 146400 79872 146405 79928
rect 146339 79867 146405 79872
rect 147254 79868 147260 79932
rect 147324 79906 147356 79932
rect 147412 79906 147417 79962
rect 151307 79962 151373 79967
rect 147324 79901 147417 79906
rect 147995 79930 148061 79933
rect 148174 79930 148180 79932
rect 147995 79928 148180 79930
rect 147324 79870 147368 79901
rect 147995 79872 148000 79928
rect 148056 79872 148180 79928
rect 147995 79870 148180 79872
rect 147324 79868 147330 79870
rect 147995 79867 148061 79870
rect 148174 79868 148180 79870
rect 148244 79868 148250 79932
rect 148731 79930 148797 79933
rect 148910 79930 148916 79932
rect 148731 79928 148916 79930
rect 148731 79872 148736 79928
rect 148792 79872 148916 79928
rect 148731 79870 148916 79872
rect 148731 79867 148797 79870
rect 148910 79868 148916 79870
rect 148980 79868 148986 79932
rect 149094 79868 149100 79932
rect 149164 79930 149170 79932
rect 149835 79930 149901 79933
rect 149164 79928 149901 79930
rect 149164 79872 149840 79928
rect 149896 79872 149901 79928
rect 149164 79870 149901 79872
rect 149164 79868 149170 79870
rect 149835 79867 149901 79870
rect 150203 79894 150269 79899
rect 145598 79732 145604 79796
rect 145668 79794 145674 79796
rect 146112 79794 146172 79867
rect 145668 79734 146172 79794
rect 145668 79732 145674 79734
rect 145465 79658 145531 79661
rect 145238 79656 145531 79658
rect 145238 79600 145470 79656
rect 145526 79600 145531 79656
rect 145238 79598 145531 79600
rect 146342 79658 146402 79867
rect 150203 79838 150208 79894
rect 150264 79838 150269 79894
rect 150382 79868 150388 79932
rect 150452 79930 150458 79932
rect 150452 79870 150510 79930
rect 150452 79868 150458 79870
rect 150750 79868 150756 79932
rect 150820 79930 150826 79932
rect 151031 79930 151097 79933
rect 151307 79932 151312 79962
rect 151368 79932 151373 79962
rect 150820 79928 151097 79930
rect 150820 79872 151036 79928
rect 151092 79872 151097 79928
rect 150820 79870 151097 79872
rect 150820 79868 150826 79870
rect 150203 79833 150269 79838
rect 150387 79838 150392 79868
rect 150448 79838 150453 79868
rect 151031 79867 151097 79870
rect 151302 79868 151308 79932
rect 151372 79930 151378 79932
rect 151494 79930 151554 80004
rect 158946 79967 159006 80142
rect 159766 80140 159772 80204
rect 159836 80140 159842 80204
rect 159774 79967 159834 80140
rect 163224 79967 163284 80278
rect 171358 80276 171364 80278
rect 171428 80276 171434 80340
rect 171542 80276 171548 80340
rect 171612 80338 171618 80340
rect 174629 80338 174695 80341
rect 171612 80336 174695 80338
rect 171612 80280 174634 80336
rect 174690 80280 174695 80336
rect 171612 80278 174695 80280
rect 171612 80276 171618 80278
rect 174629 80275 174695 80278
rect 165102 80140 165108 80204
rect 165172 80202 165178 80204
rect 171726 80202 171732 80204
rect 165172 80142 165584 80202
rect 165172 80140 165178 80142
rect 165524 79967 165584 80142
rect 169894 80142 171732 80202
rect 169518 80066 169524 80068
rect 169296 80006 169524 80066
rect 152227 79962 152293 79967
rect 151767 79930 151833 79933
rect 151372 79870 151430 79930
rect 151494 79928 151833 79930
rect 151494 79872 151772 79928
rect 151828 79872 151833 79928
rect 152227 79906 152232 79962
rect 152288 79906 152293 79962
rect 152227 79901 152293 79906
rect 152411 79962 152477 79967
rect 152411 79906 152416 79962
rect 152472 79906 152477 79962
rect 153147 79962 153213 79967
rect 152411 79901 152477 79906
rect 152595 79928 152661 79933
rect 152871 79930 152937 79933
rect 151494 79870 151833 79872
rect 151372 79868 151378 79870
rect 151767 79867 151833 79870
rect 150387 79833 150453 79838
rect 147627 79826 147693 79831
rect 147438 79732 147444 79796
rect 147508 79794 147514 79796
rect 147627 79794 147632 79826
rect 147508 79770 147632 79794
rect 147688 79770 147693 79826
rect 147508 79765 147693 79770
rect 147508 79734 147690 79765
rect 147508 79732 147514 79734
rect 148358 79732 148364 79796
rect 148428 79794 148434 79796
rect 148915 79794 148981 79797
rect 148428 79792 148981 79794
rect 148428 79736 148920 79792
rect 148976 79736 148981 79792
rect 148428 79734 148981 79736
rect 148428 79732 148434 79734
rect 148915 79731 148981 79734
rect 148961 79658 149027 79661
rect 146342 79656 149027 79658
rect 146342 79600 148966 79656
rect 149022 79600 149027 79656
rect 146342 79598 149027 79600
rect 143717 79595 143783 79598
rect 145097 79595 145163 79598
rect 145465 79595 145531 79598
rect 148961 79595 149027 79598
rect 149462 79596 149468 79660
rect 149532 79658 149538 79660
rect 150206 79658 150266 79833
rect 152230 79797 152290 79901
rect 150847 79794 150913 79797
rect 151721 79794 151787 79797
rect 150847 79792 151787 79794
rect 150847 79736 150852 79792
rect 150908 79736 151726 79792
rect 151782 79736 151787 79792
rect 150847 79734 151787 79736
rect 150847 79731 150913 79734
rect 151721 79731 151787 79734
rect 152181 79792 152290 79797
rect 152181 79736 152186 79792
rect 152242 79736 152290 79792
rect 152181 79734 152290 79736
rect 152181 79731 152247 79734
rect 149532 79598 150266 79658
rect 151997 79658 152063 79661
rect 152414 79658 152474 79901
rect 152595 79872 152600 79928
rect 152656 79872 152661 79928
rect 152595 79867 152661 79872
rect 152828 79928 152937 79930
rect 152828 79872 152876 79928
rect 152932 79872 152937 79928
rect 153147 79906 153152 79962
rect 153208 79930 153213 79962
rect 153883 79962 153949 79967
rect 153208 79906 153348 79930
rect 153147 79901 153348 79906
rect 153883 79906 153888 79962
rect 153944 79906 153949 79962
rect 154435 79962 154501 79967
rect 153883 79901 153949 79906
rect 152828 79867 152937 79872
rect 153150 79870 153348 79901
rect 152598 79797 152658 79867
rect 152598 79792 152707 79797
rect 152828 79796 152888 79867
rect 152598 79736 152646 79792
rect 152702 79736 152707 79792
rect 152598 79734 152707 79736
rect 152641 79731 152707 79734
rect 152774 79732 152780 79796
rect 152844 79734 152888 79796
rect 153009 79794 153075 79797
rect 153142 79794 153148 79796
rect 153009 79792 153148 79794
rect 153009 79736 153014 79792
rect 153070 79736 153148 79792
rect 153009 79734 153148 79736
rect 152844 79732 152850 79734
rect 153009 79731 153075 79734
rect 153142 79732 153148 79734
rect 153212 79732 153218 79796
rect 151997 79656 152474 79658
rect 151997 79600 152002 79656
rect 152058 79600 152474 79656
rect 151997 79598 152474 79600
rect 153101 79658 153167 79661
rect 153288 79658 153348 79870
rect 153886 79794 153946 79901
rect 154246 79868 154252 79932
rect 154316 79930 154322 79932
rect 154435 79930 154440 79962
rect 154316 79906 154440 79930
rect 154496 79906 154501 79962
rect 155079 79962 155145 79967
rect 154316 79901 154501 79906
rect 154316 79870 154498 79901
rect 154316 79868 154322 79870
rect 154614 79868 154620 79932
rect 154684 79930 154690 79932
rect 154895 79930 154961 79933
rect 154684 79928 154961 79930
rect 154684 79872 154900 79928
rect 154956 79872 154961 79928
rect 155079 79906 155084 79962
rect 155140 79930 155145 79962
rect 155539 79962 155605 79967
rect 155350 79930 155356 79932
rect 155140 79906 155356 79930
rect 155079 79901 155356 79906
rect 154684 79870 154961 79872
rect 155082 79870 155356 79901
rect 154684 79868 154690 79870
rect 154895 79867 154961 79870
rect 155350 79868 155356 79870
rect 155420 79868 155426 79932
rect 155539 79906 155544 79962
rect 155600 79906 155605 79962
rect 157287 79962 157353 79967
rect 155539 79901 155605 79906
rect 155723 79930 155789 79933
rect 155723 79928 155970 79930
rect 154665 79794 154731 79797
rect 153886 79792 154731 79794
rect 153886 79736 154670 79792
rect 154726 79736 154731 79792
rect 153886 79734 154731 79736
rect 154665 79731 154731 79734
rect 155033 79794 155099 79797
rect 155542 79794 155602 79901
rect 155723 79872 155728 79928
rect 155784 79872 155970 79928
rect 155723 79870 155970 79872
rect 155723 79867 155789 79870
rect 155910 79797 155970 79870
rect 156091 79928 156157 79933
rect 156091 79872 156096 79928
rect 156152 79872 156157 79928
rect 156091 79867 156157 79872
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 156643 79930 156709 79933
rect 156524 79928 156709 79930
rect 156524 79872 156648 79928
rect 156704 79872 156709 79928
rect 156524 79870 156709 79872
rect 156524 79868 156530 79870
rect 156643 79867 156709 79870
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157103 79930 157169 79933
rect 156892 79928 157169 79930
rect 156892 79872 157108 79928
rect 157164 79872 157169 79928
rect 157287 79906 157292 79962
rect 157348 79906 157353 79962
rect 158943 79962 159009 79967
rect 157287 79901 157353 79906
rect 156892 79870 157169 79872
rect 156892 79868 156898 79870
rect 157103 79867 157169 79870
rect 155033 79792 155602 79794
rect 155033 79736 155038 79792
rect 155094 79736 155602 79792
rect 155033 79734 155602 79736
rect 155861 79792 155970 79797
rect 155861 79736 155866 79792
rect 155922 79736 155970 79792
rect 155861 79734 155970 79736
rect 155033 79731 155099 79734
rect 155861 79731 155927 79734
rect 156094 79661 156154 79867
rect 156367 79794 156433 79797
rect 156367 79792 156568 79794
rect 156367 79736 156372 79792
rect 156428 79736 156568 79792
rect 156367 79734 156568 79736
rect 156367 79731 156433 79734
rect 153101 79656 153348 79658
rect 153101 79600 153106 79656
rect 153162 79600 153348 79656
rect 153101 79598 153348 79600
rect 149532 79596 149538 79598
rect 151997 79595 152063 79598
rect 153101 79595 153167 79598
rect 155534 79596 155540 79660
rect 155604 79658 155610 79660
rect 155677 79658 155743 79661
rect 155604 79656 155743 79658
rect 155604 79600 155682 79656
rect 155738 79600 155743 79656
rect 155604 79598 155743 79600
rect 155604 79596 155610 79598
rect 155677 79595 155743 79598
rect 156045 79656 156154 79661
rect 156045 79600 156050 79656
rect 156106 79600 156154 79656
rect 156045 79598 156154 79600
rect 156508 79658 156568 79734
rect 156638 79732 156644 79796
rect 156708 79794 156714 79796
rect 157290 79794 157350 79901
rect 157926 79868 157932 79932
rect 157996 79930 158002 79932
rect 158391 79930 158457 79933
rect 158575 79930 158641 79933
rect 157996 79928 158457 79930
rect 157996 79872 158396 79928
rect 158452 79872 158457 79928
rect 157996 79870 158457 79872
rect 157996 79868 158002 79870
rect 158391 79867 158457 79870
rect 158532 79928 158641 79930
rect 158532 79872 158580 79928
rect 158636 79872 158641 79928
rect 158943 79906 158948 79962
rect 159004 79906 159009 79962
rect 158943 79901 159009 79906
rect 159771 79962 159837 79967
rect 159771 79906 159776 79962
rect 159832 79906 159837 79962
rect 159771 79901 159837 79906
rect 160047 79962 160113 79967
rect 160507 79964 160573 79967
rect 160047 79906 160052 79962
rect 160108 79906 160113 79962
rect 160372 79962 160573 79964
rect 160372 79932 160512 79962
rect 160047 79901 160113 79906
rect 158532 79867 158641 79872
rect 158532 79796 158592 79867
rect 156708 79734 157350 79794
rect 156708 79732 156714 79734
rect 158478 79732 158484 79796
rect 158548 79734 158592 79796
rect 158548 79732 158554 79734
rect 158846 79732 158852 79796
rect 158916 79794 158922 79796
rect 160050 79794 160110 79901
rect 160318 79868 160324 79932
rect 160388 79906 160512 79932
rect 160568 79906 160573 79962
rect 160388 79904 160573 79906
rect 160388 79870 160432 79904
rect 160507 79901 160573 79904
rect 160875 79962 160941 79967
rect 161335 79964 161401 79967
rect 160875 79906 160880 79962
rect 160936 79906 160941 79962
rect 161292 79962 161401 79964
rect 160875 79901 160941 79906
rect 160388 79868 160394 79870
rect 158916 79734 160110 79794
rect 158916 79732 158922 79734
rect 160878 79661 160938 79901
rect 161054 79868 161060 79932
rect 161124 79930 161130 79932
rect 161292 79930 161340 79962
rect 161124 79906 161340 79930
rect 161396 79906 161401 79962
rect 161124 79901 161401 79906
rect 161519 79964 161585 79967
rect 162991 79964 163057 79967
rect 161519 79962 161858 79964
rect 161519 79906 161524 79962
rect 161580 79932 161858 79962
rect 162948 79962 163057 79964
rect 161979 79932 162045 79933
rect 161580 79906 161796 79932
rect 161519 79904 161796 79906
rect 161519 79901 161585 79904
rect 161124 79870 161352 79901
rect 161124 79868 161130 79870
rect 161790 79868 161796 79904
rect 161860 79868 161866 79932
rect 161974 79868 161980 79932
rect 162044 79930 162050 79932
rect 162044 79870 162136 79930
rect 162044 79868 162050 79870
rect 162342 79868 162348 79932
rect 162412 79930 162418 79932
rect 162623 79930 162689 79933
rect 162412 79928 162689 79930
rect 162412 79872 162628 79928
rect 162684 79872 162689 79928
rect 162412 79870 162689 79872
rect 162412 79868 162418 79870
rect 161979 79867 162045 79868
rect 162623 79867 162689 79870
rect 162948 79906 162996 79962
rect 163052 79906 163057 79962
rect 162948 79901 163057 79906
rect 163175 79962 163284 79967
rect 163543 79964 163609 79967
rect 163175 79906 163180 79962
rect 163236 79906 163284 79962
rect 163500 79962 163609 79964
rect 163500 79932 163548 79962
rect 163175 79904 163284 79906
rect 163175 79901 163241 79904
rect 162948 79797 163008 79901
rect 163446 79868 163452 79932
rect 163516 79906 163548 79932
rect 163604 79906 163609 79962
rect 164003 79962 164069 79967
rect 163516 79901 163609 79906
rect 163819 79930 163885 79933
rect 163819 79928 163928 79930
rect 163516 79870 163560 79901
rect 163819 79872 163824 79928
rect 163880 79872 163928 79928
rect 164003 79906 164008 79962
rect 164064 79906 164069 79962
rect 164555 79962 164621 79967
rect 164279 79930 164345 79933
rect 164555 79932 164560 79962
rect 164616 79932 164621 79962
rect 165291 79962 165357 79967
rect 165291 79932 165296 79962
rect 165352 79932 165357 79962
rect 165524 79962 165633 79967
rect 164003 79901 164069 79906
rect 164236 79928 164345 79930
rect 163516 79868 163522 79870
rect 163819 79867 163928 79872
rect 163868 79797 163928 79867
rect 161289 79794 161355 79797
rect 162393 79794 162459 79797
rect 161289 79792 162459 79794
rect 161289 79736 161294 79792
rect 161350 79736 162398 79792
rect 162454 79736 162459 79792
rect 161289 79734 162459 79736
rect 161289 79731 161355 79734
rect 162393 79731 162459 79734
rect 162715 79792 162781 79797
rect 162715 79736 162720 79792
rect 162776 79736 162781 79792
rect 162715 79731 162781 79736
rect 162945 79792 163011 79797
rect 163359 79794 163425 79797
rect 162945 79736 162950 79792
rect 163006 79736 163011 79792
rect 162945 79731 163011 79736
rect 163316 79792 163425 79794
rect 163316 79736 163364 79792
rect 163420 79736 163425 79792
rect 163316 79731 163425 79736
rect 163865 79792 163931 79797
rect 163865 79736 163870 79792
rect 163926 79736 163931 79792
rect 163865 79731 163931 79736
rect 156781 79658 156847 79661
rect 156508 79656 156847 79658
rect 156508 79600 156786 79656
rect 156842 79600 156847 79656
rect 156508 79598 156847 79600
rect 160878 79656 160987 79661
rect 160878 79600 160926 79656
rect 160982 79600 160987 79656
rect 160878 79598 160987 79600
rect 156045 79595 156111 79598
rect 156781 79595 156847 79598
rect 160921 79595 160987 79598
rect 161381 79658 161447 79661
rect 161841 79658 161907 79661
rect 161381 79656 161907 79658
rect 161381 79600 161386 79656
rect 161442 79600 161846 79656
rect 161902 79600 161907 79656
rect 161381 79598 161907 79600
rect 161381 79595 161447 79598
rect 161841 79595 161907 79598
rect 162526 79596 162532 79660
rect 162596 79658 162602 79660
rect 162718 79658 162778 79731
rect 163316 79660 163376 79731
rect 162596 79598 162778 79658
rect 162596 79596 162602 79598
rect 163262 79596 163268 79660
rect 163332 79598 163376 79660
rect 163332 79596 163338 79598
rect 163446 79596 163452 79660
rect 163516 79658 163522 79660
rect 164006 79658 164066 79901
rect 164236 79872 164284 79928
rect 164340 79872 164345 79928
rect 164236 79867 164345 79872
rect 164550 79868 164556 79932
rect 164620 79930 164626 79932
rect 164620 79870 164678 79930
rect 164620 79868 164626 79870
rect 165286 79868 165292 79932
rect 165356 79930 165362 79932
rect 165356 79870 165414 79930
rect 165524 79906 165572 79962
rect 165628 79906 165633 79962
rect 168787 79962 168853 79967
rect 165524 79904 165633 79906
rect 165567 79901 165633 79904
rect 166671 79930 166737 79933
rect 167315 79932 167381 79933
rect 167683 79932 167749 79933
rect 167867 79932 167933 79933
rect 166942 79930 166948 79932
rect 166671 79928 166948 79930
rect 166671 79872 166676 79928
rect 166732 79872 166948 79928
rect 166671 79870 166948 79872
rect 165356 79868 165362 79870
rect 166671 79867 166737 79870
rect 166942 79868 166948 79870
rect 167012 79868 167018 79932
rect 167310 79930 167316 79932
rect 167224 79870 167316 79930
rect 167310 79868 167316 79870
rect 167380 79868 167386 79932
rect 167678 79930 167684 79932
rect 167592 79870 167684 79930
rect 167678 79868 167684 79870
rect 167748 79868 167754 79932
rect 167862 79868 167868 79932
rect 167932 79930 167938 79932
rect 167932 79870 168024 79930
rect 168235 79928 168301 79933
rect 168419 79932 168485 79933
rect 168787 79932 168792 79962
rect 168848 79932 168853 79962
rect 168235 79872 168240 79928
rect 168296 79872 168301 79928
rect 167932 79868 167938 79870
rect 167315 79867 167381 79868
rect 167683 79867 167749 79868
rect 167867 79867 167933 79868
rect 168235 79867 168301 79872
rect 168414 79868 168420 79932
rect 168484 79930 168490 79932
rect 168484 79870 168576 79930
rect 168484 79868 168490 79870
rect 168782 79868 168788 79932
rect 168852 79930 168858 79932
rect 168971 79930 169037 79933
rect 169150 79930 169156 79932
rect 168852 79870 168910 79930
rect 168971 79928 169156 79930
rect 168971 79872 168976 79928
rect 169032 79872 169156 79928
rect 168971 79870 169156 79872
rect 168852 79868 168858 79870
rect 168419 79867 168485 79868
rect 168971 79867 169037 79870
rect 169150 79868 169156 79870
rect 169220 79868 169226 79932
rect 169296 79930 169356 80006
rect 169518 80004 169524 80006
rect 169588 80004 169594 80068
rect 169894 79967 169954 80142
rect 171726 80140 171732 80142
rect 171796 80140 171802 80204
rect 178309 80202 178375 80205
rect 172470 80200 178375 80202
rect 172470 80144 178314 80200
rect 178370 80144 178375 80200
rect 172470 80142 178375 80144
rect 170806 80066 170812 80068
rect 170446 80006 170812 80066
rect 169891 79962 169957 79967
rect 169431 79930 169497 79933
rect 169296 79928 169497 79930
rect 169296 79872 169436 79928
rect 169492 79872 169497 79928
rect 169296 79870 169497 79872
rect 169431 79867 169497 79870
rect 169615 79928 169681 79933
rect 169615 79872 169620 79928
rect 169676 79872 169681 79928
rect 169891 79906 169896 79962
rect 169952 79906 169957 79962
rect 170075 79962 170141 79967
rect 170075 79932 170080 79962
rect 170136 79932 170141 79962
rect 170446 79933 170506 80006
rect 170806 80004 170812 80006
rect 170876 80004 170882 80068
rect 172470 80066 172530 80142
rect 178309 80139 178375 80142
rect 171504 80006 172530 80066
rect 171504 79967 171564 80006
rect 172830 80004 172836 80068
rect 172900 80004 172906 80068
rect 173014 80004 173020 80068
rect 173084 80066 173090 80068
rect 173084 80006 173496 80066
rect 173084 80004 173090 80006
rect 171455 79962 171564 79967
rect 169891 79901 169957 79906
rect 169615 79867 169681 79872
rect 170070 79868 170076 79932
rect 170140 79930 170146 79932
rect 170140 79870 170198 79930
rect 170259 79928 170325 79933
rect 170259 79872 170264 79928
rect 170320 79872 170325 79928
rect 170140 79868 170146 79870
rect 170259 79867 170325 79872
rect 170443 79928 170509 79933
rect 170719 79930 170785 79933
rect 170443 79872 170448 79928
rect 170504 79872 170509 79928
rect 170443 79867 170509 79872
rect 170676 79928 170785 79930
rect 170676 79872 170724 79928
rect 170780 79872 170785 79928
rect 170676 79867 170785 79872
rect 170903 79930 170969 79933
rect 171179 79932 171245 79933
rect 170903 79928 171104 79930
rect 170903 79872 170908 79928
rect 170964 79872 171104 79928
rect 170903 79870 171104 79872
rect 170903 79867 170969 79870
rect 164236 79794 164296 79867
rect 164236 79734 165400 79794
rect 165340 79661 165400 79734
rect 165654 79732 165660 79796
rect 165724 79794 165730 79796
rect 166211 79794 166277 79797
rect 165724 79792 166277 79794
rect 165724 79736 166216 79792
rect 166272 79736 166277 79792
rect 165724 79734 166277 79736
rect 165724 79732 165730 79734
rect 166211 79731 166277 79734
rect 166395 79792 166461 79797
rect 166395 79736 166400 79792
rect 166456 79736 166461 79792
rect 166395 79731 166461 79736
rect 168046 79732 168052 79796
rect 168116 79794 168122 79796
rect 168238 79794 168298 79867
rect 168116 79734 168298 79794
rect 168557 79794 168623 79797
rect 168833 79794 168899 79797
rect 168557 79792 168899 79794
rect 168557 79736 168562 79792
rect 168618 79736 168838 79792
rect 168894 79736 168899 79792
rect 168557 79734 168899 79736
rect 168116 79732 168122 79734
rect 168557 79731 168623 79734
rect 168833 79731 168899 79734
rect 169017 79792 169083 79797
rect 169017 79736 169022 79792
rect 169078 79736 169083 79792
rect 169017 79731 169083 79736
rect 169618 79794 169678 79867
rect 169886 79794 169892 79796
rect 169618 79734 169892 79794
rect 169886 79732 169892 79734
rect 169956 79732 169962 79796
rect 164233 79660 164299 79661
rect 163516 79598 164066 79658
rect 163516 79596 163522 79598
rect 164182 79596 164188 79660
rect 164252 79658 164299 79660
rect 164252 79656 164344 79658
rect 164294 79600 164344 79656
rect 164252 79598 164344 79600
rect 165337 79656 165403 79661
rect 165337 79600 165342 79656
rect 165398 79600 165403 79656
rect 164252 79596 164299 79598
rect 164233 79595 164299 79596
rect 165337 79595 165403 79600
rect 165705 79658 165771 79661
rect 165838 79658 165844 79660
rect 165705 79656 165844 79658
rect 165705 79600 165710 79656
rect 165766 79600 165844 79656
rect 165705 79598 165844 79600
rect 165705 79595 165771 79598
rect 165838 79596 165844 79598
rect 165908 79596 165914 79660
rect 166257 79658 166323 79661
rect 166398 79658 166458 79731
rect 166257 79656 166458 79658
rect 166257 79600 166262 79656
rect 166318 79600 166458 79656
rect 166257 79598 166458 79600
rect 166257 79595 166323 79598
rect 166758 79596 166764 79660
rect 166828 79658 166834 79660
rect 166901 79658 166967 79661
rect 166828 79656 166967 79658
rect 166828 79600 166906 79656
rect 166962 79600 166967 79656
rect 166828 79598 166967 79600
rect 169020 79658 169080 79731
rect 170262 79661 170322 79867
rect 170121 79658 170187 79661
rect 169020 79656 170187 79658
rect 169020 79600 170126 79656
rect 170182 79600 170187 79656
rect 169020 79598 170187 79600
rect 170262 79656 170371 79661
rect 170489 79660 170555 79661
rect 170262 79600 170310 79656
rect 170366 79600 170371 79656
rect 170262 79598 170371 79600
rect 166828 79596 166834 79598
rect 166901 79595 166967 79598
rect 170121 79595 170187 79598
rect 170305 79595 170371 79598
rect 170438 79596 170444 79660
rect 170508 79658 170555 79660
rect 170676 79658 170736 79867
rect 171044 79796 171104 79870
rect 171174 79868 171180 79932
rect 171244 79930 171250 79932
rect 171244 79870 171336 79930
rect 171455 79906 171460 79962
rect 171516 79906 171564 79962
rect 171455 79904 171564 79906
rect 171639 79930 171705 79933
rect 172283 79932 172349 79933
rect 172467 79932 172533 79933
rect 171910 79930 171916 79932
rect 171639 79928 171916 79930
rect 171455 79901 171521 79904
rect 171639 79872 171644 79928
rect 171700 79872 171916 79928
rect 171639 79870 171916 79872
rect 171244 79868 171250 79870
rect 171179 79867 171245 79868
rect 171639 79867 171705 79870
rect 171910 79868 171916 79870
rect 171980 79868 171986 79932
rect 172278 79930 172284 79932
rect 172192 79870 172284 79930
rect 172278 79868 172284 79870
rect 172348 79868 172354 79932
rect 172462 79868 172468 79932
rect 172532 79930 172538 79932
rect 172838 79930 172898 80004
rect 173295 79930 173361 79933
rect 172532 79870 172624 79930
rect 172838 79928 173361 79930
rect 172838 79872 173300 79928
rect 173356 79872 173361 79928
rect 172838 79870 173361 79872
rect 172532 79868 172538 79870
rect 172283 79867 172349 79868
rect 172467 79867 172533 79868
rect 173295 79867 173361 79870
rect 170990 79732 170996 79796
rect 171060 79734 171104 79796
rect 171593 79794 171659 79797
rect 172094 79794 172100 79796
rect 171593 79792 172100 79794
rect 171593 79736 171598 79792
rect 171654 79736 172100 79792
rect 171593 79734 172100 79736
rect 171060 79732 171066 79734
rect 171593 79731 171659 79734
rect 172094 79732 172100 79734
rect 172164 79732 172170 79796
rect 172462 79732 172468 79796
rect 172532 79794 172538 79796
rect 172743 79794 172809 79797
rect 172532 79792 172809 79794
rect 172532 79736 172748 79792
rect 172804 79736 172809 79792
rect 172532 79734 172809 79736
rect 173436 79794 173496 80006
rect 173755 79930 173821 79933
rect 173755 79928 174186 79930
rect 173755 79872 173760 79928
rect 173816 79872 174186 79928
rect 173755 79870 174186 79872
rect 173755 79867 173821 79870
rect 173663 79794 173729 79797
rect 173436 79792 173729 79794
rect 173436 79736 173668 79792
rect 173724 79736 173729 79792
rect 173436 79734 173729 79736
rect 174126 79794 174186 79870
rect 174261 79794 174327 79797
rect 174126 79792 174327 79794
rect 174126 79736 174266 79792
rect 174322 79736 174327 79792
rect 174126 79734 174327 79736
rect 172532 79732 172538 79734
rect 172743 79731 172809 79734
rect 173663 79731 173729 79734
rect 174261 79731 174327 79734
rect 171041 79658 171107 79661
rect 170508 79656 170600 79658
rect 170550 79600 170600 79656
rect 170508 79598 170600 79600
rect 170676 79656 171107 79658
rect 170676 79600 171046 79656
rect 171102 79600 171107 79656
rect 170676 79598 171107 79600
rect 170508 79596 170555 79598
rect 170489 79595 170555 79596
rect 171041 79595 171107 79598
rect 171501 79658 171567 79661
rect 178493 79658 178559 79661
rect 171501 79656 178559 79658
rect 171501 79600 171506 79656
rect 171562 79600 178498 79656
rect 178554 79600 178559 79656
rect 171501 79598 178559 79600
rect 171501 79595 171567 79598
rect 178493 79595 178559 79598
rect 6913 79522 6979 79525
rect 172973 79522 173039 79525
rect 6913 79520 173039 79522
rect 6913 79464 6918 79520
rect 6974 79464 172978 79520
rect 173034 79464 173039 79520
rect 6913 79462 173039 79464
rect 6913 79459 6979 79462
rect 172973 79459 173039 79462
rect 3785 79386 3851 79389
rect 174537 79386 174603 79389
rect 3785 79384 174603 79386
rect 3785 79328 3790 79384
rect 3846 79328 174542 79384
rect 174598 79328 174603 79384
rect 3785 79326 174603 79328
rect 3785 79323 3851 79326
rect 174537 79323 174603 79326
rect 3601 79250 3667 79253
rect 173341 79250 173407 79253
rect 3601 79248 173407 79250
rect 3601 79192 3606 79248
rect 3662 79192 173346 79248
rect 173402 79192 173407 79248
rect 3601 79190 173407 79192
rect 3601 79187 3667 79190
rect 173341 79187 173407 79190
rect 3417 79114 3483 79117
rect 173249 79114 173315 79117
rect 3417 79112 173315 79114
rect 3417 79056 3422 79112
rect 3478 79056 173254 79112
rect 173310 79056 173315 79112
rect 3417 79054 173315 79056
rect 3417 79051 3483 79054
rect 173249 79051 173315 79054
rect 173382 79052 173388 79116
rect 173452 79114 173458 79116
rect 173525 79114 173591 79117
rect 173452 79112 173591 79114
rect 173452 79056 173530 79112
rect 173586 79056 173591 79112
rect 173452 79054 173591 79056
rect 173452 79052 173458 79054
rect 173525 79051 173591 79054
rect 3233 78978 3299 78981
rect 173065 78978 173131 78981
rect 3233 78976 173131 78978
rect 3233 78920 3238 78976
rect 3294 78920 173070 78976
rect 173126 78920 173131 78976
rect 3233 78918 173131 78920
rect 3233 78915 3299 78918
rect 173065 78915 173131 78918
rect 173198 78916 173204 78980
rect 173268 78978 173274 78980
rect 173268 78918 180810 78978
rect 173268 78916 173274 78918
rect 138422 78780 138428 78844
rect 138492 78842 138498 78844
rect 138565 78842 138631 78845
rect 145925 78844 145991 78845
rect 145925 78842 145972 78844
rect 138492 78840 138631 78842
rect 138492 78784 138570 78840
rect 138626 78784 138631 78840
rect 138492 78782 138631 78784
rect 145880 78840 145972 78842
rect 145880 78784 145930 78840
rect 145880 78782 145972 78784
rect 138492 78780 138498 78782
rect 138565 78779 138631 78782
rect 145925 78780 145972 78782
rect 146036 78780 146042 78844
rect 148542 78780 148548 78844
rect 148612 78842 148618 78844
rect 149053 78842 149119 78845
rect 148612 78840 149119 78842
rect 148612 78784 149058 78840
rect 149114 78784 149119 78840
rect 148612 78782 149119 78784
rect 148612 78780 148618 78782
rect 145925 78779 145991 78780
rect 149053 78779 149119 78782
rect 149697 78842 149763 78845
rect 151353 78844 151419 78845
rect 150382 78842 150388 78844
rect 149697 78840 150388 78842
rect 149697 78784 149702 78840
rect 149758 78784 150388 78840
rect 149697 78782 150388 78784
rect 149697 78779 149763 78782
rect 150382 78780 150388 78782
rect 150452 78780 150458 78844
rect 151302 78780 151308 78844
rect 151372 78842 151419 78844
rect 157241 78842 157307 78845
rect 163497 78842 163563 78845
rect 151372 78840 151464 78842
rect 151414 78784 151464 78840
rect 151372 78782 151464 78784
rect 157241 78840 163563 78842
rect 157241 78784 157246 78840
rect 157302 78784 163502 78840
rect 163558 78784 163563 78840
rect 157241 78782 163563 78784
rect 151372 78780 151419 78782
rect 151353 78779 151419 78780
rect 157241 78779 157307 78782
rect 163497 78779 163563 78782
rect 165429 78844 165495 78845
rect 165429 78840 165476 78844
rect 165540 78842 165546 78844
rect 165429 78784 165434 78840
rect 165429 78780 165476 78784
rect 165540 78782 165586 78842
rect 165540 78780 165546 78782
rect 168414 78780 168420 78844
rect 168484 78842 168490 78844
rect 172094 78842 172100 78844
rect 168484 78782 172100 78842
rect 168484 78780 168490 78782
rect 172094 78780 172100 78782
rect 172164 78780 172170 78844
rect 180750 78842 180810 78918
rect 397453 78842 397519 78845
rect 180750 78840 397519 78842
rect 180750 78784 397458 78840
rect 397514 78784 397519 78840
rect 180750 78782 397519 78784
rect 165429 78779 165495 78780
rect 397453 78779 397519 78782
rect 144310 78644 144316 78708
rect 144380 78706 144386 78708
rect 144637 78706 144703 78709
rect 144380 78704 144703 78706
rect 144380 78648 144642 78704
rect 144698 78648 144703 78704
rect 144380 78646 144703 78648
rect 144380 78644 144386 78646
rect 144637 78643 144703 78646
rect 145230 78644 145236 78708
rect 145300 78706 145306 78708
rect 146201 78706 146267 78709
rect 145300 78704 146267 78706
rect 145300 78648 146206 78704
rect 146262 78648 146267 78704
rect 145300 78646 146267 78648
rect 145300 78644 145306 78646
rect 146201 78643 146267 78646
rect 147070 78644 147076 78708
rect 147140 78706 147146 78708
rect 147397 78706 147463 78709
rect 148777 78708 148843 78709
rect 148726 78706 148732 78708
rect 147140 78704 147463 78706
rect 147140 78648 147402 78704
rect 147458 78648 147463 78704
rect 147140 78646 147463 78648
rect 148686 78646 148732 78706
rect 148796 78704 148843 78708
rect 149053 78708 149119 78709
rect 149053 78706 149100 78708
rect 148838 78648 148843 78704
rect 147140 78644 147146 78646
rect 147397 78643 147463 78646
rect 148726 78644 148732 78646
rect 148796 78644 148843 78648
rect 149008 78704 149100 78706
rect 149008 78648 149058 78704
rect 149008 78646 149100 78648
rect 148777 78643 148843 78644
rect 149053 78644 149100 78646
rect 149164 78644 149170 78708
rect 149646 78644 149652 78708
rect 149716 78706 149722 78708
rect 150249 78706 150315 78709
rect 149716 78704 150315 78706
rect 149716 78648 150254 78704
rect 150310 78648 150315 78704
rect 149716 78646 150315 78648
rect 149716 78644 149722 78646
rect 149053 78643 149119 78644
rect 150249 78643 150315 78646
rect 150433 78706 150499 78709
rect 150750 78706 150756 78708
rect 150433 78704 150756 78706
rect 150433 78648 150438 78704
rect 150494 78648 150756 78704
rect 150433 78646 150756 78648
rect 150433 78643 150499 78646
rect 150750 78644 150756 78646
rect 150820 78644 150826 78708
rect 151169 78706 151235 78709
rect 151670 78706 151676 78708
rect 151169 78704 151676 78706
rect 151169 78648 151174 78704
rect 151230 78648 151676 78704
rect 151169 78646 151676 78648
rect 151169 78643 151235 78646
rect 151670 78644 151676 78646
rect 151740 78644 151746 78708
rect 153878 78644 153884 78708
rect 153948 78706 153954 78708
rect 154205 78706 154271 78709
rect 153948 78704 154271 78706
rect 153948 78648 154210 78704
rect 154266 78648 154271 78704
rect 153948 78646 154271 78648
rect 153948 78644 153954 78646
rect 154205 78643 154271 78646
rect 159030 78644 159036 78708
rect 159100 78706 159106 78708
rect 159725 78706 159791 78709
rect 160277 78708 160343 78709
rect 160277 78706 160324 78708
rect 159100 78704 159791 78706
rect 159100 78648 159730 78704
rect 159786 78648 159791 78704
rect 159100 78646 159791 78648
rect 160232 78704 160324 78706
rect 160232 78648 160282 78704
rect 160232 78646 160324 78648
rect 159100 78644 159106 78646
rect 159725 78643 159791 78646
rect 160277 78644 160324 78646
rect 160388 78644 160394 78708
rect 161013 78706 161079 78709
rect 161238 78706 161244 78708
rect 161013 78704 161244 78706
rect 161013 78648 161018 78704
rect 161074 78648 161244 78704
rect 161013 78646 161244 78648
rect 160277 78643 160343 78644
rect 161013 78643 161079 78646
rect 161238 78644 161244 78646
rect 161308 78644 161314 78708
rect 161565 78706 161631 78709
rect 161790 78706 161796 78708
rect 161565 78704 161796 78706
rect 161565 78648 161570 78704
rect 161626 78648 161796 78704
rect 161565 78646 161796 78648
rect 161565 78643 161631 78646
rect 161790 78644 161796 78646
rect 161860 78644 161866 78708
rect 162158 78644 162164 78708
rect 162228 78706 162234 78708
rect 162485 78706 162551 78709
rect 162228 78704 162551 78706
rect 162228 78648 162490 78704
rect 162546 78648 162551 78704
rect 162228 78646 162551 78648
rect 162228 78644 162234 78646
rect 162485 78643 162551 78646
rect 162669 78708 162735 78709
rect 162669 78704 162716 78708
rect 162780 78706 162786 78708
rect 163221 78706 163287 78709
rect 164785 78706 164851 78709
rect 165613 78708 165679 78709
rect 165797 78708 165863 78709
rect 165613 78706 165660 78708
rect 162669 78648 162674 78704
rect 162669 78644 162716 78648
rect 162780 78646 162826 78706
rect 163221 78704 164851 78706
rect 163221 78648 163226 78704
rect 163282 78648 164790 78704
rect 164846 78648 164851 78704
rect 163221 78646 164851 78648
rect 165568 78704 165660 78706
rect 165568 78648 165618 78704
rect 165568 78646 165660 78648
rect 162780 78644 162786 78646
rect 162669 78643 162735 78644
rect 163221 78643 163287 78646
rect 164785 78643 164851 78646
rect 165613 78644 165660 78646
rect 165724 78644 165730 78708
rect 165797 78704 165844 78708
rect 165908 78706 165914 78708
rect 165797 78648 165802 78704
rect 165797 78644 165844 78648
rect 165908 78646 165954 78706
rect 165908 78644 165914 78646
rect 166390 78644 166396 78708
rect 166460 78706 166466 78708
rect 166717 78706 166783 78709
rect 166460 78704 166783 78706
rect 166460 78648 166722 78704
rect 166778 78648 166783 78704
rect 166460 78646 166783 78648
rect 166460 78644 166466 78646
rect 165613 78643 165679 78644
rect 165797 78643 165863 78644
rect 166717 78643 166783 78646
rect 167678 78644 167684 78708
rect 167748 78706 167754 78708
rect 168005 78706 168071 78709
rect 167748 78704 168071 78706
rect 167748 78648 168010 78704
rect 168066 78648 168071 78704
rect 167748 78646 168071 78648
rect 167748 78644 167754 78646
rect 168005 78643 168071 78646
rect 169845 78706 169911 78709
rect 170070 78706 170076 78708
rect 169845 78704 170076 78706
rect 169845 78648 169850 78704
rect 169906 78648 170076 78704
rect 169845 78646 170076 78648
rect 169845 78643 169911 78646
rect 170070 78644 170076 78646
rect 170140 78644 170146 78708
rect 170438 78644 170444 78708
rect 170508 78706 170514 78708
rect 170581 78706 170647 78709
rect 170508 78704 170647 78706
rect 170508 78648 170586 78704
rect 170642 78648 170647 78704
rect 170508 78646 170647 78648
rect 170508 78644 170514 78646
rect 170581 78643 170647 78646
rect 170857 78706 170923 78709
rect 171542 78706 171548 78708
rect 170857 78704 171548 78706
rect 170857 78648 170862 78704
rect 170918 78648 171548 78704
rect 170857 78646 171548 78648
rect 170857 78643 170923 78646
rect 171542 78644 171548 78646
rect 171612 78644 171618 78708
rect 171777 78706 171843 78709
rect 172145 78706 172211 78709
rect 171777 78704 172211 78706
rect 171777 78648 171782 78704
rect 171838 78648 172150 78704
rect 172206 78648 172211 78704
rect 171777 78646 172211 78648
rect 171777 78643 171843 78646
rect 172145 78643 172211 78646
rect 172329 78706 172395 78709
rect 462313 78706 462379 78709
rect 172329 78704 462379 78706
rect 172329 78648 172334 78704
rect 172390 78648 462318 78704
rect 462374 78648 462379 78704
rect 172329 78646 462379 78648
rect 172329 78643 172395 78646
rect 462313 78643 462379 78646
rect 145414 78508 145420 78572
rect 145484 78570 145490 78572
rect 146109 78570 146175 78573
rect 145484 78568 146175 78570
rect 145484 78512 146114 78568
rect 146170 78512 146175 78568
rect 145484 78510 146175 78512
rect 145484 78508 145490 78510
rect 146109 78507 146175 78510
rect 149830 78508 149836 78572
rect 149900 78570 149906 78572
rect 150157 78570 150223 78573
rect 149900 78568 150223 78570
rect 149900 78512 150162 78568
rect 150218 78512 150223 78568
rect 149900 78510 150223 78512
rect 149900 78508 149906 78510
rect 150157 78507 150223 78510
rect 151302 78508 151308 78572
rect 151372 78570 151378 78572
rect 151721 78570 151787 78573
rect 151372 78568 151787 78570
rect 151372 78512 151726 78568
rect 151782 78512 151787 78568
rect 151372 78510 151787 78512
rect 151372 78508 151378 78510
rect 151721 78507 151787 78510
rect 158662 78508 158668 78572
rect 158732 78570 158738 78572
rect 158805 78570 158871 78573
rect 158732 78568 158871 78570
rect 158732 78512 158810 78568
rect 158866 78512 158871 78568
rect 158732 78510 158871 78512
rect 158732 78508 158738 78510
rect 158805 78507 158871 78510
rect 161054 78508 161060 78572
rect 161124 78570 161130 78572
rect 161197 78570 161263 78573
rect 161124 78568 161263 78570
rect 161124 78512 161202 78568
rect 161258 78512 161263 78568
rect 161124 78510 161263 78512
rect 161124 78508 161130 78510
rect 161197 78507 161263 78510
rect 164918 78508 164924 78572
rect 164988 78570 164994 78572
rect 165521 78570 165587 78573
rect 164988 78568 165587 78570
rect 164988 78512 165526 78568
rect 165582 78512 165587 78568
rect 164988 78510 165587 78512
rect 164988 78508 164994 78510
rect 165521 78507 165587 78510
rect 167637 78570 167703 78573
rect 169569 78572 169635 78573
rect 167862 78570 167868 78572
rect 167637 78568 167868 78570
rect 167637 78512 167642 78568
rect 167698 78512 167868 78568
rect 167637 78510 167868 78512
rect 167637 78507 167703 78510
rect 167862 78508 167868 78510
rect 167932 78508 167938 78572
rect 169518 78508 169524 78572
rect 169588 78570 169635 78572
rect 170857 78570 170923 78573
rect 170990 78570 170996 78572
rect 169588 78568 169680 78570
rect 169630 78512 169680 78568
rect 169588 78510 169680 78512
rect 170857 78568 170996 78570
rect 170857 78512 170862 78568
rect 170918 78512 170996 78568
rect 170857 78510 170996 78512
rect 169588 78508 169635 78510
rect 169569 78507 169635 78508
rect 170857 78507 170923 78510
rect 170990 78508 170996 78510
rect 171060 78508 171066 78572
rect 172237 78570 172303 78573
rect 396717 78570 396783 78573
rect 172237 78568 396783 78570
rect 172237 78512 172242 78568
rect 172298 78512 396722 78568
rect 396778 78512 396783 78568
rect 172237 78510 396783 78512
rect 172237 78507 172303 78510
rect 396717 78507 396783 78510
rect 148869 78434 148935 78437
rect 150014 78434 150020 78436
rect 148869 78432 150020 78434
rect 148869 78376 148874 78432
rect 148930 78376 150020 78432
rect 148869 78374 150020 78376
rect 148869 78371 148935 78374
rect 150014 78372 150020 78374
rect 150084 78372 150090 78436
rect 160870 78372 160876 78436
rect 160940 78434 160946 78436
rect 161473 78434 161539 78437
rect 160940 78432 161539 78434
rect 160940 78376 161478 78432
rect 161534 78376 161539 78432
rect 160940 78374 161539 78376
rect 160940 78372 160946 78374
rect 161473 78371 161539 78374
rect 162117 78434 162183 78437
rect 168741 78434 168807 78437
rect 162117 78432 168807 78434
rect 162117 78376 162122 78432
rect 162178 78376 168746 78432
rect 168802 78376 168807 78432
rect 162117 78374 168807 78376
rect 162117 78371 162183 78374
rect 168741 78371 168807 78374
rect 171501 78434 171567 78437
rect 172697 78434 172763 78437
rect 396574 78434 396580 78436
rect 171501 78432 172530 78434
rect 171501 78376 171506 78432
rect 171562 78376 172530 78432
rect 171501 78374 172530 78376
rect 171501 78371 171567 78374
rect 157149 78298 157215 78301
rect 172329 78298 172395 78301
rect 157149 78296 172395 78298
rect 157149 78240 157154 78296
rect 157210 78240 172334 78296
rect 172390 78240 172395 78296
rect 157149 78238 172395 78240
rect 172470 78298 172530 78374
rect 172697 78432 396580 78434
rect 172697 78376 172702 78432
rect 172758 78376 396580 78432
rect 172697 78374 396580 78376
rect 172697 78371 172763 78374
rect 396574 78372 396580 78374
rect 396644 78372 396650 78436
rect 173985 78298 174051 78301
rect 172470 78296 174051 78298
rect 172470 78240 173990 78296
rect 174046 78240 174051 78296
rect 172470 78238 174051 78240
rect 157149 78235 157215 78238
rect 172329 78235 172395 78238
rect 173985 78235 174051 78238
rect 127985 78162 128051 78165
rect 130009 78164 130075 78165
rect 128670 78162 128676 78164
rect 127985 78160 128676 78162
rect 127985 78104 127990 78160
rect 128046 78104 128676 78160
rect 127985 78102 128676 78104
rect 127985 78099 128051 78102
rect 128670 78100 128676 78102
rect 128740 78100 128746 78164
rect 129958 78162 129964 78164
rect 129918 78102 129964 78162
rect 130028 78160 130075 78164
rect 130070 78104 130075 78160
rect 129958 78100 129964 78102
rect 130028 78100 130075 78104
rect 130009 78099 130075 78100
rect 137829 78164 137895 78165
rect 137829 78160 137876 78164
rect 137940 78162 137946 78164
rect 155033 78162 155099 78165
rect 155350 78162 155356 78164
rect 137829 78104 137834 78160
rect 137829 78100 137876 78104
rect 137940 78102 137986 78162
rect 155033 78160 155356 78162
rect 155033 78104 155038 78160
rect 155094 78104 155356 78160
rect 155033 78102 155356 78104
rect 137940 78100 137946 78102
rect 137829 78099 137895 78100
rect 155033 78099 155099 78102
rect 155350 78100 155356 78102
rect 155420 78100 155426 78164
rect 158294 78100 158300 78164
rect 158364 78162 158370 78164
rect 158529 78162 158595 78165
rect 158364 78160 158595 78162
rect 158364 78104 158534 78160
rect 158590 78104 158595 78160
rect 158364 78102 158595 78104
rect 158364 78100 158370 78102
rect 158529 78099 158595 78102
rect 159766 78100 159772 78164
rect 159836 78162 159842 78164
rect 166625 78162 166691 78165
rect 159836 78160 166691 78162
rect 159836 78104 166630 78160
rect 166686 78104 166691 78160
rect 159836 78102 166691 78104
rect 159836 78100 159842 78102
rect 166625 78099 166691 78102
rect 167085 78162 167151 78165
rect 167310 78162 167316 78164
rect 167085 78160 167316 78162
rect 167085 78104 167090 78160
rect 167146 78104 167316 78160
rect 167085 78102 167316 78104
rect 167085 78099 167151 78102
rect 167310 78100 167316 78102
rect 167380 78100 167386 78164
rect 167678 78100 167684 78164
rect 167748 78162 167754 78164
rect 168189 78162 168255 78165
rect 167748 78160 168255 78162
rect 167748 78104 168194 78160
rect 168250 78104 168255 78160
rect 167748 78102 168255 78104
rect 167748 78100 167754 78102
rect 168189 78099 168255 78102
rect 168649 78162 168715 78165
rect 168782 78162 168788 78164
rect 168649 78160 168788 78162
rect 168649 78104 168654 78160
rect 168710 78104 168788 78160
rect 168649 78102 168788 78104
rect 168649 78099 168715 78102
rect 168782 78100 168788 78102
rect 168852 78100 168858 78164
rect 168925 78162 168991 78165
rect 169150 78162 169156 78164
rect 168925 78160 169156 78162
rect 168925 78104 168930 78160
rect 168986 78104 169156 78160
rect 168925 78102 169156 78104
rect 168925 78099 168991 78102
rect 169150 78100 169156 78102
rect 169220 78100 169226 78164
rect 169518 78100 169524 78164
rect 169588 78162 169594 78164
rect 169661 78162 169727 78165
rect 169588 78160 169727 78162
rect 169588 78104 169666 78160
rect 169722 78104 169727 78160
rect 169588 78102 169727 78104
rect 169588 78100 169594 78102
rect 169661 78099 169727 78102
rect 170213 78162 170279 78165
rect 172237 78162 172303 78165
rect 170213 78160 172303 78162
rect 170213 78104 170218 78160
rect 170274 78104 172242 78160
rect 172298 78104 172303 78160
rect 170213 78102 172303 78104
rect 170213 78099 170279 78102
rect 172237 78099 172303 78102
rect 128721 78028 128787 78029
rect 128670 78026 128676 78028
rect 128630 77966 128676 78026
rect 128740 78024 128787 78028
rect 128782 77968 128787 78024
rect 128670 77964 128676 77966
rect 128740 77964 128787 77968
rect 128721 77963 128787 77964
rect 129733 78028 129799 78029
rect 130101 78028 130167 78029
rect 130469 78028 130535 78029
rect 131021 78028 131087 78029
rect 129733 78024 129780 78028
rect 129844 78026 129850 78028
rect 129733 77968 129738 78024
rect 129733 77964 129780 77968
rect 129844 77966 129890 78026
rect 130101 78024 130148 78028
rect 130212 78026 130218 78028
rect 130469 78026 130516 78028
rect 130101 77968 130106 78024
rect 129844 77964 129850 77966
rect 130101 77964 130148 77968
rect 130212 77966 130258 78026
rect 130424 78024 130516 78026
rect 130424 77968 130474 78024
rect 130424 77966 130516 77968
rect 130212 77964 130218 77966
rect 130469 77964 130516 77966
rect 130580 77964 130586 78028
rect 131021 78024 131068 78028
rect 131132 78026 131138 78028
rect 135529 78026 135595 78029
rect 135662 78026 135668 78028
rect 131021 77968 131026 78024
rect 131021 77964 131068 77968
rect 131132 77966 131178 78026
rect 135529 78024 135668 78026
rect 135529 77968 135534 78024
rect 135590 77968 135668 78024
rect 135529 77966 135668 77968
rect 131132 77964 131138 77966
rect 129733 77963 129799 77964
rect 130101 77963 130167 77964
rect 130469 77963 130535 77964
rect 131021 77963 131087 77964
rect 135529 77963 135595 77966
rect 135662 77964 135668 77966
rect 135732 77964 135738 78028
rect 136398 77964 136404 78028
rect 136468 78026 136474 78028
rect 138013 78026 138079 78029
rect 136468 78024 138079 78026
rect 136468 77968 138018 78024
rect 138074 77968 138079 78024
rect 136468 77966 138079 77968
rect 136468 77964 136474 77966
rect 138013 77963 138079 77966
rect 158110 77964 158116 78028
rect 158180 78026 158186 78028
rect 158437 78026 158503 78029
rect 158180 78024 158503 78026
rect 158180 77968 158442 78024
rect 158498 77968 158503 78024
rect 158180 77966 158503 77968
rect 158180 77964 158186 77966
rect 158437 77963 158503 77966
rect 159173 78026 159239 78029
rect 161197 78026 161263 78029
rect 159173 78024 161263 78026
rect 159173 77968 159178 78024
rect 159234 77968 161202 78024
rect 161258 77968 161263 78024
rect 159173 77966 161263 77968
rect 159173 77963 159239 77966
rect 161197 77963 161263 77966
rect 162853 78026 162919 78029
rect 478873 78026 478939 78029
rect 162853 78024 478939 78026
rect 162853 77968 162858 78024
rect 162914 77968 478878 78024
rect 478934 77968 478939 78024
rect 162853 77966 478939 77968
rect 162853 77963 162919 77966
rect 478873 77963 478939 77966
rect 150985 77890 151051 77893
rect 137970 77888 151051 77890
rect 137970 77832 150990 77888
rect 151046 77832 151051 77888
rect 137970 77830 151051 77832
rect 137970 77754 138030 77830
rect 150985 77827 151051 77830
rect 156413 77890 156479 77893
rect 170213 77890 170279 77893
rect 156413 77888 170279 77890
rect 156413 77832 156418 77888
rect 156474 77832 170218 77888
rect 170274 77832 170279 77888
rect 156413 77830 170279 77832
rect 156413 77827 156479 77830
rect 170213 77827 170279 77830
rect 171358 77828 171364 77892
rect 171428 77890 171434 77892
rect 483013 77890 483079 77893
rect 171428 77888 483079 77890
rect 171428 77832 483018 77888
rect 483074 77832 483079 77888
rect 171428 77830 483079 77832
rect 171428 77828 171434 77830
rect 483013 77827 483079 77830
rect 133462 77694 138030 77754
rect 131982 77556 131988 77620
rect 132052 77618 132058 77620
rect 133462 77618 133522 77694
rect 163078 77692 163084 77756
rect 163148 77754 163154 77756
rect 163589 77754 163655 77757
rect 163148 77752 163655 77754
rect 163148 77696 163594 77752
rect 163650 77696 163655 77752
rect 163148 77694 163655 77696
rect 163148 77692 163154 77694
rect 163589 77691 163655 77694
rect 166625 77754 166691 77757
rect 166625 77752 168482 77754
rect 166625 77696 166630 77752
rect 166686 77696 168482 77752
rect 166625 77694 168482 77696
rect 166625 77691 166691 77694
rect 132052 77558 133522 77618
rect 163129 77618 163195 77621
rect 163262 77618 163268 77620
rect 163129 77616 163268 77618
rect 163129 77560 163134 77616
rect 163190 77560 163268 77616
rect 163129 77558 163268 77560
rect 132052 77556 132058 77558
rect 163129 77555 163195 77558
rect 163262 77556 163268 77558
rect 163332 77556 163338 77620
rect 164550 77556 164556 77620
rect 164620 77618 164626 77620
rect 165061 77618 165127 77621
rect 166809 77620 166875 77621
rect 168097 77620 168163 77621
rect 166758 77618 166764 77620
rect 164620 77616 165127 77618
rect 164620 77560 165066 77616
rect 165122 77560 165127 77616
rect 164620 77558 165127 77560
rect 166718 77558 166764 77618
rect 166828 77616 166875 77620
rect 168046 77618 168052 77620
rect 166870 77560 166875 77616
rect 164620 77556 164626 77558
rect 165061 77555 165127 77558
rect 166758 77556 166764 77558
rect 166828 77556 166875 77560
rect 168006 77558 168052 77618
rect 168116 77616 168163 77620
rect 168158 77560 168163 77616
rect 168046 77556 168052 77558
rect 168116 77556 168163 77560
rect 168422 77618 168482 77694
rect 168422 77558 170322 77618
rect 166809 77555 166875 77556
rect 168097 77555 168163 77556
rect 132861 77482 132927 77485
rect 133086 77482 133092 77484
rect 132861 77480 133092 77482
rect 132861 77424 132866 77480
rect 132922 77424 133092 77480
rect 132861 77422 133092 77424
rect 132861 77419 132927 77422
rect 133086 77420 133092 77422
rect 133156 77420 133162 77484
rect 148174 77420 148180 77484
rect 148244 77482 148250 77484
rect 148869 77482 148935 77485
rect 157057 77484 157123 77485
rect 157006 77482 157012 77484
rect 148244 77480 148935 77482
rect 148244 77424 148874 77480
rect 148930 77424 148935 77480
rect 148244 77422 148935 77424
rect 156966 77422 157012 77482
rect 157076 77480 157123 77484
rect 157118 77424 157123 77480
rect 148244 77420 148250 77422
rect 148869 77419 148935 77422
rect 157006 77420 157012 77422
rect 157076 77420 157123 77424
rect 157057 77419 157123 77420
rect 152590 77284 152596 77348
rect 152660 77346 152666 77348
rect 153009 77346 153075 77349
rect 152660 77344 153075 77346
rect 152660 77288 153014 77344
rect 153070 77288 153075 77344
rect 152660 77286 153075 77288
rect 152660 77284 152666 77286
rect 153009 77283 153075 77286
rect 161974 77148 161980 77212
rect 162044 77210 162050 77212
rect 162209 77210 162275 77213
rect 162044 77208 162275 77210
rect 162044 77152 162214 77208
rect 162270 77152 162275 77208
rect 162044 77150 162275 77152
rect 170262 77210 170322 77558
rect 171961 77346 172027 77349
rect 170814 77344 172027 77346
rect 170814 77288 171966 77344
rect 172022 77288 172027 77344
rect 170814 77286 172027 77288
rect 170814 77210 170874 77286
rect 171961 77283 172027 77286
rect 172278 77284 172284 77348
rect 172348 77346 172354 77348
rect 178769 77346 178835 77349
rect 172348 77344 178835 77346
rect 172348 77288 178774 77344
rect 178830 77288 178835 77344
rect 172348 77286 178835 77288
rect 172348 77284 172354 77286
rect 178769 77283 178835 77286
rect 170262 77150 170874 77210
rect 171869 77210 171935 77213
rect 172462 77210 172468 77212
rect 171869 77208 172468 77210
rect 171869 77152 171874 77208
rect 171930 77152 172468 77208
rect 171869 77150 172468 77152
rect 162044 77148 162050 77150
rect 162209 77147 162275 77150
rect 171869 77147 171935 77150
rect 172462 77148 172468 77150
rect 172532 77148 172538 77212
rect 142470 77012 142476 77076
rect 142540 77074 142546 77076
rect 170213 77074 170279 77077
rect 142540 77072 170279 77074
rect 142540 77016 170218 77072
rect 170274 77016 170279 77072
rect 142540 77014 170279 77016
rect 142540 77012 142546 77014
rect 170213 77011 170279 77014
rect 111793 76938 111859 76941
rect 134149 76938 134215 76941
rect 111793 76936 134215 76938
rect 111793 76880 111798 76936
rect 111854 76880 134154 76936
rect 134210 76880 134215 76936
rect 111793 76878 134215 76880
rect 111793 76875 111859 76878
rect 134149 76875 134215 76878
rect 144729 76938 144795 76941
rect 247033 76938 247099 76941
rect 144729 76936 247099 76938
rect 144729 76880 144734 76936
rect 144790 76880 247038 76936
rect 247094 76880 247099 76936
rect 144729 76878 247099 76880
rect 144729 76875 144795 76878
rect 247033 76875 247099 76878
rect 93853 76802 93919 76805
rect 132585 76802 132651 76805
rect 93853 76800 132651 76802
rect 93853 76744 93858 76800
rect 93914 76744 132590 76800
rect 132646 76744 132651 76800
rect 93853 76742 132651 76744
rect 93853 76739 93919 76742
rect 132585 76739 132651 76742
rect 147673 76802 147739 76805
rect 282913 76802 282979 76805
rect 147673 76800 282979 76802
rect 147673 76744 147678 76800
rect 147734 76744 282918 76800
rect 282974 76744 282979 76800
rect 147673 76742 282979 76744
rect 147673 76739 147739 76742
rect 282913 76739 282979 76742
rect 20713 76666 20779 76669
rect 127249 76666 127315 76669
rect 20713 76664 127315 76666
rect 20713 76608 20718 76664
rect 20774 76608 127254 76664
rect 127310 76608 127315 76664
rect 20713 76606 127315 76608
rect 20713 76603 20779 76606
rect 127249 76603 127315 76606
rect 152825 76666 152891 76669
rect 152958 76666 152964 76668
rect 152825 76664 152964 76666
rect 152825 76608 152830 76664
rect 152886 76608 152964 76664
rect 152825 76606 152964 76608
rect 152825 76603 152891 76606
rect 152958 76604 152964 76606
rect 153028 76604 153034 76668
rect 170213 76666 170279 76669
rect 173249 76666 173315 76669
rect 549253 76666 549319 76669
rect 170213 76664 173315 76666
rect 170213 76608 170218 76664
rect 170274 76608 173254 76664
rect 173310 76608 173315 76664
rect 170213 76606 173315 76608
rect 170213 76603 170279 76606
rect 173249 76603 173315 76606
rect 173390 76664 549319 76666
rect 173390 76608 549258 76664
rect 549314 76608 549319 76664
rect 173390 76606 549319 76608
rect 1393 76530 1459 76533
rect 125685 76530 125751 76533
rect 1393 76528 125751 76530
rect 1393 76472 1398 76528
rect 1454 76472 125690 76528
rect 125746 76472 125751 76528
rect 1393 76470 125751 76472
rect 1393 76467 1459 76470
rect 125685 76467 125751 76470
rect 128353 76530 128419 76533
rect 128854 76530 128860 76532
rect 128353 76528 128860 76530
rect 128353 76472 128358 76528
rect 128414 76472 128860 76528
rect 128353 76470 128860 76472
rect 128353 76467 128419 76470
rect 128854 76468 128860 76470
rect 128924 76468 128930 76532
rect 168833 76530 168899 76533
rect 173390 76530 173450 76606
rect 549253 76603 549319 76606
rect 565813 76530 565879 76533
rect 168833 76528 173450 76530
rect 168833 76472 168838 76528
rect 168894 76472 173450 76528
rect 168833 76470 173450 76472
rect 176610 76528 565879 76530
rect 176610 76472 565818 76528
rect 565874 76472 565879 76528
rect 176610 76470 565879 76472
rect 168833 76467 168899 76470
rect 169886 76332 169892 76396
rect 169956 76394 169962 76396
rect 176610 76394 176670 76470
rect 565813 76467 565879 76470
rect 169956 76334 176670 76394
rect 169956 76332 169962 76334
rect 155718 76196 155724 76260
rect 155788 76258 155794 76260
rect 155861 76258 155927 76261
rect 155788 76256 155927 76258
rect 155788 76200 155866 76256
rect 155922 76200 155927 76256
rect 155788 76198 155927 76200
rect 155788 76196 155794 76198
rect 155861 76195 155927 76198
rect 142613 76122 142679 76125
rect 142838 76122 142844 76124
rect 142613 76120 142844 76122
rect 142613 76064 142618 76120
rect 142674 76064 142844 76120
rect 142613 76062 142844 76064
rect 142613 76059 142679 76062
rect 142838 76060 142844 76062
rect 142908 76060 142914 76124
rect 125777 75988 125843 75989
rect 125726 75986 125732 75988
rect 125686 75926 125732 75986
rect 125796 75984 125843 75988
rect 125838 75928 125843 75984
rect 125726 75924 125732 75926
rect 125796 75924 125843 75928
rect 140262 75924 140268 75988
rect 140332 75986 140338 75988
rect 140589 75986 140655 75989
rect 140332 75984 140655 75986
rect 140332 75928 140594 75984
rect 140650 75928 140655 75984
rect 140332 75926 140655 75928
rect 140332 75924 140338 75926
rect 125777 75923 125843 75924
rect 140589 75923 140655 75926
rect 142838 75924 142844 75988
rect 142908 75986 142914 75988
rect 143257 75986 143323 75989
rect 143809 75988 143875 75989
rect 142908 75984 143323 75986
rect 142908 75928 143262 75984
rect 143318 75928 143323 75984
rect 142908 75926 143323 75928
rect 142908 75924 142914 75926
rect 143257 75923 143323 75926
rect 143758 75924 143764 75988
rect 143828 75986 143875 75988
rect 154389 75988 154455 75989
rect 143828 75984 143920 75986
rect 143870 75928 143920 75984
rect 143828 75926 143920 75928
rect 154389 75984 154436 75988
rect 154500 75986 154506 75988
rect 154389 75928 154394 75984
rect 143828 75924 143875 75926
rect 143809 75923 143875 75924
rect 154389 75924 154436 75928
rect 154500 75926 154546 75986
rect 154500 75924 154506 75926
rect 154614 75924 154620 75988
rect 154684 75986 154690 75988
rect 155217 75986 155283 75989
rect 154684 75984 155283 75986
rect 154684 75928 155222 75984
rect 155278 75928 155283 75984
rect 154684 75926 155283 75928
rect 154684 75924 154690 75926
rect 154389 75923 154455 75924
rect 155217 75923 155283 75926
rect 156137 75986 156203 75989
rect 156454 75986 156460 75988
rect 156137 75984 156460 75986
rect 156137 75928 156142 75984
rect 156198 75928 156460 75984
rect 156137 75926 156460 75928
rect 156137 75923 156203 75926
rect 156454 75924 156460 75926
rect 156524 75924 156530 75988
rect 171133 75986 171199 75989
rect 171910 75986 171916 75988
rect 171133 75984 171916 75986
rect 171133 75928 171138 75984
rect 171194 75928 171916 75984
rect 171133 75926 171916 75928
rect 171133 75923 171199 75926
rect 171910 75924 171916 75926
rect 171980 75924 171986 75988
rect 140078 75788 140084 75852
rect 140148 75850 140154 75852
rect 140405 75850 140471 75853
rect 140148 75848 140471 75850
rect 140148 75792 140410 75848
rect 140466 75792 140471 75848
rect 140148 75790 140471 75792
rect 140148 75788 140154 75790
rect 140405 75787 140471 75790
rect 154062 75788 154068 75852
rect 154132 75850 154138 75852
rect 154481 75850 154547 75853
rect 154132 75848 154547 75850
rect 154132 75792 154486 75848
rect 154542 75792 154547 75848
rect 154132 75790 154547 75792
rect 154132 75788 154138 75790
rect 154481 75787 154547 75790
rect 139117 75714 139183 75717
rect 173893 75714 173959 75717
rect 139117 75712 173959 75714
rect 139117 75656 139122 75712
rect 139178 75656 173898 75712
rect 173954 75656 173959 75712
rect 139117 75654 173959 75656
rect 139117 75651 139183 75654
rect 173893 75651 173959 75654
rect 57973 75578 58039 75581
rect 130326 75578 130332 75580
rect 57973 75576 130332 75578
rect 57973 75520 57978 75576
rect 58034 75520 130332 75576
rect 57973 75518 130332 75520
rect 57973 75515 58039 75518
rect 130326 75516 130332 75518
rect 130396 75516 130402 75580
rect 139945 75578 140011 75581
rect 176653 75578 176719 75581
rect 139945 75576 176719 75578
rect 139945 75520 139950 75576
rect 140006 75520 176658 75576
rect 176714 75520 176719 75576
rect 139945 75518 176719 75520
rect 139945 75515 140011 75518
rect 176653 75515 176719 75518
rect 53833 75442 53899 75445
rect 129774 75442 129780 75444
rect 53833 75440 129780 75442
rect 53833 75384 53838 75440
rect 53894 75384 129780 75440
rect 53833 75382 129780 75384
rect 53833 75379 53899 75382
rect 129774 75380 129780 75382
rect 129844 75380 129850 75444
rect 156873 75442 156939 75445
rect 402973 75442 403039 75445
rect 156873 75440 403039 75442
rect 156873 75384 156878 75440
rect 156934 75384 402978 75440
rect 403034 75384 403039 75440
rect 156873 75382 403039 75384
rect 156873 75379 156939 75382
rect 402973 75379 403039 75382
rect 35893 75306 35959 75309
rect 123661 75306 123727 75309
rect 35893 75304 123727 75306
rect 35893 75248 35898 75304
rect 35954 75248 123666 75304
rect 123722 75248 123727 75304
rect 35893 75246 123727 75248
rect 35893 75243 35959 75246
rect 123661 75243 123727 75246
rect 164141 75306 164207 75309
rect 496813 75306 496879 75309
rect 164141 75304 496879 75306
rect 164141 75248 164146 75304
rect 164202 75248 496818 75304
rect 496874 75248 496879 75304
rect 164141 75246 496879 75248
rect 164141 75243 164207 75246
rect 496813 75243 496879 75246
rect 2773 75170 2839 75173
rect 125542 75170 125548 75172
rect 2773 75168 125548 75170
rect 2773 75112 2778 75168
rect 2834 75112 125548 75168
rect 2773 75110 125548 75112
rect 2773 75107 2839 75110
rect 125542 75108 125548 75110
rect 125612 75108 125618 75172
rect 167126 75108 167132 75172
rect 167196 75170 167202 75172
rect 528553 75170 528619 75173
rect 167196 75168 528619 75170
rect 167196 75112 528558 75168
rect 528614 75112 528619 75168
rect 167196 75110 528619 75112
rect 167196 75108 167202 75110
rect 528553 75107 528619 75110
rect 130377 74490 130443 74493
rect 135294 74490 135300 74492
rect 130377 74488 135300 74490
rect 130377 74432 130382 74488
rect 130438 74432 135300 74488
rect 130377 74430 135300 74432
rect 130377 74427 130443 74430
rect 135294 74428 135300 74430
rect 135364 74428 135370 74492
rect 140681 74082 140747 74085
rect 194593 74082 194659 74085
rect 140681 74080 194659 74082
rect 140681 74024 140686 74080
rect 140742 74024 194598 74080
rect 194654 74024 194659 74080
rect 140681 74022 194659 74024
rect 140681 74019 140747 74022
rect 194593 74019 194659 74022
rect 144126 73884 144132 73948
rect 144196 73946 144202 73948
rect 230473 73946 230539 73949
rect 144196 73944 230539 73946
rect 144196 73888 230478 73944
rect 230534 73888 230539 73944
rect 144196 73886 230539 73888
rect 144196 73884 144202 73886
rect 230473 73883 230539 73886
rect 40033 73810 40099 73813
rect 127985 73810 128051 73813
rect 40033 73808 128051 73810
rect 40033 73752 40038 73808
rect 40094 73752 127990 73808
rect 128046 73752 128051 73808
rect 40033 73750 128051 73752
rect 40033 73747 40099 73750
rect 127985 73747 128051 73750
rect 144678 73748 144684 73812
rect 144748 73810 144754 73812
rect 244273 73810 244339 73813
rect 144748 73808 244339 73810
rect 144748 73752 244278 73808
rect 244334 73752 244339 73808
rect 144748 73750 244339 73752
rect 144748 73748 144754 73750
rect 244273 73747 244339 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 162158 72660 162164 72724
rect 162228 72722 162234 72724
rect 178677 72722 178743 72725
rect 162228 72720 178743 72722
rect 162228 72664 178682 72720
rect 178738 72664 178743 72720
rect 162228 72662 178743 72664
rect 162228 72660 162234 72662
rect 178677 72659 178743 72662
rect 147438 72524 147444 72588
rect 147508 72586 147514 72588
rect 284293 72586 284359 72589
rect 147508 72584 284359 72586
rect 147508 72528 284298 72584
rect 284354 72528 284359 72584
rect 147508 72526 284359 72528
rect 147508 72524 147514 72526
rect 284293 72523 284359 72526
rect 148910 72388 148916 72452
rect 148980 72450 148986 72452
rect 298093 72450 298159 72453
rect 148980 72448 298159 72450
rect 148980 72392 298098 72448
rect 298154 72392 298159 72448
rect 148980 72390 298159 72392
rect 148980 72388 148986 72390
rect 298093 72387 298159 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 153142 71164 153148 71228
rect 153212 71226 153218 71228
rect 353293 71226 353359 71229
rect 153212 71224 353359 71226
rect 153212 71168 353298 71224
rect 353354 71168 353359 71224
rect 153212 71166 353359 71168
rect 153212 71164 153218 71166
rect 353293 71163 353359 71166
rect 163446 71028 163452 71092
rect 163516 71090 163522 71092
rect 494053 71090 494119 71093
rect 163516 71088 494119 71090
rect 163516 71032 494058 71088
rect 494114 71032 494119 71088
rect 163516 71030 494119 71032
rect 163516 71028 163522 71030
rect 494053 71027 494119 71030
rect 138974 69532 138980 69596
rect 139044 69594 139050 69596
rect 175273 69594 175339 69597
rect 139044 69592 175339 69594
rect 139044 69536 175278 69592
rect 175334 69536 175339 69592
rect 139044 69534 175339 69536
rect 139044 69532 139050 69534
rect 175273 69531 175339 69534
rect 165470 68172 165476 68236
rect 165540 68234 165546 68236
rect 511993 68234 512059 68237
rect 165540 68232 512059 68234
rect 165540 68176 511998 68232
rect 512054 68176 512059 68232
rect 165540 68174 512059 68176
rect 165540 68172 165546 68174
rect 511993 68171 512059 68174
rect 140262 65452 140268 65516
rect 140332 65514 140338 65516
rect 193213 65514 193279 65517
rect 140332 65512 193279 65514
rect 140332 65456 193218 65512
rect 193274 65456 193279 65512
rect 140332 65454 193279 65456
rect 140332 65452 140338 65454
rect 193213 65451 193279 65454
rect 166390 62868 166396 62932
rect 166460 62930 166466 62932
rect 529933 62930 529999 62933
rect 166460 62928 529999 62930
rect 166460 62872 529938 62928
rect 529994 62872 529999 62928
rect 166460 62870 529999 62872
rect 166460 62868 166466 62870
rect 529933 62867 529999 62870
rect 172094 62732 172100 62796
rect 172164 62794 172170 62796
rect 550633 62794 550699 62797
rect 172164 62792 550699 62794
rect 172164 62736 550638 62792
rect 550694 62736 550699 62792
rect 172164 62734 550699 62736
rect 172164 62732 172170 62734
rect 550633 62731 550699 62734
rect 160686 61372 160692 61436
rect 160756 61434 160762 61436
rect 459553 61434 459619 61437
rect 160756 61432 459619 61434
rect 160756 61376 459558 61432
rect 459614 61376 459619 61432
rect 160756 61374 459619 61376
rect 160756 61372 160762 61374
rect 459553 61371 459619 61374
rect 138606 60012 138612 60076
rect 138676 60074 138682 60076
rect 172513 60074 172579 60077
rect 138676 60072 172579 60074
rect 138676 60016 172518 60072
rect 172574 60016 172579 60072
rect 138676 60014 172579 60016
rect 138676 60012 138682 60014
rect 172513 60011 172579 60014
rect 143022 59876 143028 59940
rect 143092 59938 143098 59940
rect 227713 59938 227779 59941
rect 143092 59936 227779 59938
rect 143092 59880 227718 59936
rect 227774 59880 227779 59936
rect 143092 59878 227779 59880
rect 143092 59876 143098 59878
rect 227713 59875 227779 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 149462 53076 149468 53140
rect 149532 53138 149538 53140
rect 316033 53138 316099 53141
rect 149532 53136 316099 53138
rect 149532 53080 316038 53136
rect 316094 53080 316099 53136
rect 149532 53078 316099 53080
rect 149532 53076 149538 53078
rect 316033 53075 316099 53078
rect 152590 47500 152596 47564
rect 152660 47562 152666 47564
rect 351913 47562 351979 47565
rect 152660 47560 351979 47562
rect 152660 47504 351918 47560
rect 351974 47504 351979 47560
rect 152660 47502 351979 47504
rect 152660 47500 152666 47502
rect 351913 47499 351979 47502
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 127065 44978 127131 44981
rect 135662 44978 135668 44980
rect 127065 44976 135668 44978
rect 127065 44920 127070 44976
rect 127126 44920 135668 44976
rect 127065 44918 135668 44920
rect 127065 44915 127131 44918
rect 135662 44916 135668 44918
rect 135732 44916 135738 44980
rect 91093 44842 91159 44845
rect 133270 44842 133276 44844
rect 91093 44840 133276 44842
rect 91093 44784 91098 44840
rect 91154 44784 133276 44840
rect 91093 44782 133276 44784
rect 91093 44779 91159 44782
rect 133270 44780 133276 44782
rect 133340 44780 133346 44844
rect 147254 44780 147260 44844
rect 147324 44842 147330 44844
rect 280153 44842 280219 44845
rect 147324 44840 280219 44842
rect 147324 44784 280158 44840
rect 280214 44784 280219 44840
rect 147324 44782 280219 44784
rect 147324 44780 147330 44782
rect 280153 44779 280219 44782
rect 22093 43482 22159 43485
rect 127198 43482 127204 43484
rect 22093 43480 127204 43482
rect 22093 43424 22098 43480
rect 22154 43424 127204 43480
rect 22093 43422 127204 43424
rect 22093 43419 22159 43422
rect 127198 43420 127204 43422
rect 127268 43420 127274 43484
rect 153878 40564 153884 40628
rect 153948 40626 153954 40628
rect 367093 40626 367159 40629
rect 153948 40624 367159 40626
rect 153948 40568 367098 40624
rect 367154 40568 367159 40624
rect 153948 40566 367159 40568
rect 153948 40564 153954 40566
rect 367093 40563 367159 40566
rect 154062 35124 154068 35188
rect 154132 35186 154138 35188
rect 372613 35186 372679 35189
rect 154132 35184 372679 35186
rect 154132 35128 372618 35184
rect 372674 35128 372679 35184
rect 154132 35126 372679 35128
rect 154132 35124 154138 35126
rect 372613 35123 372679 35126
rect 143206 34036 143212 34100
rect 143276 34098 143282 34100
rect 226425 34098 226491 34101
rect 143276 34096 226491 34098
rect 143276 34040 226430 34096
rect 226486 34040 226491 34096
rect 143276 34038 226491 34040
rect 143276 34036 143282 34038
rect 226425 34035 226491 34038
rect 145230 33900 145236 33964
rect 145300 33962 145306 33964
rect 266353 33962 266419 33965
rect 145300 33960 266419 33962
rect 145300 33904 266358 33960
rect 266414 33904 266419 33960
rect 145300 33902 266419 33904
rect 145300 33900 145306 33902
rect 266353 33899 266419 33902
rect 170622 33764 170628 33828
rect 170692 33826 170698 33828
rect 578233 33826 578299 33829
rect 170692 33824 578299 33826
rect 170692 33768 578238 33824
rect 578294 33768 578299 33824
rect 170692 33766 578299 33768
rect 170692 33764 170698 33766
rect 578233 33763 578299 33766
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 166574 32540 166580 32604
rect 166644 32602 166650 32604
rect 531313 32602 531379 32605
rect 166644 32600 531379 32602
rect 166644 32544 531318 32600
rect 531374 32544 531379 32600
rect 166644 32542 531379 32544
rect 166644 32540 166650 32542
rect 531313 32539 531379 32542
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 169518 32404 169524 32468
rect 169588 32466 169594 32468
rect 567193 32466 567259 32469
rect 169588 32464 567259 32466
rect 169588 32408 567198 32464
rect 567254 32408 567259 32464
rect 169588 32406 567259 32408
rect 169588 32404 169594 32406
rect 567193 32403 567259 32406
rect 167678 30908 167684 30972
rect 167748 30970 167754 30972
rect 546493 30970 546559 30973
rect 167748 30968 546559 30970
rect 167748 30912 546498 30968
rect 546554 30912 546559 30968
rect 167748 30910 546559 30912
rect 167748 30908 167754 30910
rect 546493 30907 546559 30910
rect 149646 29548 149652 29612
rect 149716 29610 149722 29612
rect 317413 29610 317479 29613
rect 149716 29608 317479 29610
rect 149716 29552 317418 29608
rect 317474 29552 317479 29608
rect 149716 29550 317479 29552
rect 149716 29548 149722 29550
rect 317413 29547 317479 29550
rect 140446 28460 140452 28524
rect 140516 28522 140522 28524
rect 193305 28522 193371 28525
rect 140516 28520 193371 28522
rect 140516 28464 193310 28520
rect 193366 28464 193371 28520
rect 140516 28462 193371 28464
rect 140516 28460 140522 28462
rect 193305 28459 193371 28462
rect 142838 28324 142844 28388
rect 142908 28386 142914 28388
rect 229093 28386 229159 28389
rect 142908 28384 229159 28386
rect 142908 28328 229098 28384
rect 229154 28328 229159 28384
rect 142908 28326 229159 28328
rect 142908 28324 142914 28326
rect 229093 28323 229159 28326
rect 165102 28188 165108 28252
rect 165172 28250 165178 28252
rect 514845 28250 514911 28253
rect 165172 28248 514911 28250
rect 165172 28192 514850 28248
rect 514906 28192 514911 28248
rect 165172 28190 514911 28192
rect 165172 28188 165178 28190
rect 514845 28187 514911 28190
rect 165286 26964 165292 27028
rect 165356 27026 165362 27028
rect 510613 27026 510679 27029
rect 165356 27024 510679 27026
rect 165356 26968 510618 27024
rect 510674 26968 510679 27024
rect 165356 26966 510679 26968
rect 165356 26964 165362 26966
rect 510613 26963 510679 26966
rect 170806 26828 170812 26892
rect 170876 26890 170882 26892
rect 576853 26890 576919 26893
rect 170876 26888 576919 26890
rect 170876 26832 576858 26888
rect 576914 26832 576919 26888
rect 170876 26830 576919 26832
rect 170876 26828 170882 26830
rect 576853 26827 576919 26830
rect 155534 25468 155540 25532
rect 155604 25530 155610 25532
rect 386413 25530 386479 25533
rect 155604 25528 386479 25530
rect 155604 25472 386418 25528
rect 386474 25472 386479 25528
rect 155604 25470 386479 25472
rect 155604 25468 155610 25470
rect 386413 25467 386479 25470
rect 157926 24108 157932 24172
rect 157996 24170 158002 24172
rect 422293 24170 422359 24173
rect 157996 24168 422359 24170
rect 157996 24112 422298 24168
rect 422354 24112 422359 24168
rect 157996 24110 422359 24112
rect 157996 24108 158002 24110
rect 422293 24107 422359 24110
rect 170438 21660 170444 21724
rect 170508 21722 170514 21724
rect 319437 21722 319503 21725
rect 170508 21720 319503 21722
rect 170508 21664 319442 21720
rect 319498 21664 319503 21720
rect 170508 21662 319503 21664
rect 170508 21660 170514 21662
rect 319437 21659 319503 21662
rect 158846 21524 158852 21588
rect 158916 21586 158922 21588
rect 442993 21586 443059 21589
rect 158916 21584 443059 21586
rect 158916 21528 442998 21584
rect 443054 21528 443059 21584
rect 158916 21526 443059 21528
rect 158916 21524 158922 21526
rect 442993 21523 443059 21526
rect 160870 21388 160876 21452
rect 160940 21450 160946 21452
rect 460933 21450 460999 21453
rect 160940 21448 460999 21450
rect 160940 21392 460938 21448
rect 460994 21392 460999 21448
rect 160940 21390 460999 21392
rect 160940 21388 160946 21390
rect 460933 21387 460999 21390
rect 162342 21252 162348 21316
rect 162412 21314 162418 21316
rect 476113 21314 476179 21317
rect 162412 21312 476179 21314
rect 162412 21256 476118 21312
rect 476174 21256 476179 21312
rect 162412 21254 476179 21256
rect 162412 21252 162418 21254
rect 476113 21251 476179 21254
rect 144494 20164 144500 20228
rect 144564 20226 144570 20228
rect 248413 20226 248479 20229
rect 144564 20224 248479 20226
rect 144564 20168 248418 20224
rect 248474 20168 248479 20224
rect 144564 20166 248479 20168
rect 144564 20164 144570 20166
rect 248413 20163 248479 20166
rect 161054 20028 161060 20092
rect 161124 20090 161130 20092
rect 458173 20090 458239 20093
rect 161124 20088 458239 20090
rect 161124 20032 458178 20088
rect 458234 20032 458239 20088
rect 161124 20030 458239 20032
rect 161124 20028 161130 20030
rect 458173 20027 458239 20030
rect 137686 19892 137692 19956
rect 137756 19954 137762 19956
rect 160553 19954 160619 19957
rect 137756 19952 160619 19954
rect 137756 19896 160558 19952
rect 160614 19896 160619 19952
rect 137756 19894 160619 19896
rect 137756 19892 137762 19894
rect 160553 19891 160619 19894
rect 163630 19892 163636 19956
rect 163700 19954 163706 19956
rect 495433 19954 495499 19957
rect 163700 19952 495499 19954
rect 163700 19896 495438 19952
rect 495494 19896 495499 19952
rect 163700 19894 495499 19896
rect 163700 19892 163706 19894
rect 495433 19891 495499 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 4061 19410 4127 19413
rect -960 19408 4127 19410
rect -960 19352 4066 19408
rect 4122 19352 4127 19408
rect -960 19350 4127 19352
rect -960 19260 480 19350
rect 4061 19347 4127 19350
rect 140078 18940 140084 19004
rect 140148 19002 140154 19004
rect 191833 19002 191899 19005
rect 140148 19000 191899 19002
rect 140148 18944 191838 19000
rect 191894 18944 191899 19000
rect 140148 18942 191899 18944
rect 140148 18940 140154 18942
rect 191833 18939 191899 18942
rect 152774 18804 152780 18868
rect 152844 18866 152850 18868
rect 350533 18866 350599 18869
rect 152844 18864 350599 18866
rect 152844 18808 350538 18864
rect 350594 18808 350599 18864
rect 152844 18806 350599 18808
rect 152844 18804 152850 18806
rect 350533 18803 350599 18806
rect 158110 18668 158116 18732
rect 158180 18730 158186 18732
rect 423673 18730 423739 18733
rect 158180 18728 423739 18730
rect 158180 18672 423678 18728
rect 423734 18672 423739 18728
rect 158180 18670 423739 18672
rect 158180 18668 158186 18670
rect 423673 18667 423739 18670
rect 167862 18532 167868 18596
rect 167932 18594 167938 18596
rect 547873 18594 547939 18597
rect 167932 18592 547939 18594
rect 167932 18536 547878 18592
rect 547934 18536 547939 18592
rect 167932 18534 547939 18536
rect 167932 18532 167938 18534
rect 547873 18531 547939 18534
rect 156822 17308 156828 17372
rect 156892 17370 156898 17372
rect 405733 17370 405799 17373
rect 156892 17368 405799 17370
rect 156892 17312 405738 17368
rect 405794 17312 405799 17368
rect 156892 17310 405799 17312
rect 156892 17308 156898 17310
rect 405733 17307 405799 17310
rect 161238 17172 161244 17236
rect 161308 17234 161314 17236
rect 456885 17234 456951 17237
rect 161308 17232 456951 17234
rect 161308 17176 456890 17232
rect 456946 17176 456951 17232
rect 161308 17174 456951 17176
rect 161308 17172 161314 17174
rect 456885 17171 456951 17174
rect 149830 16220 149836 16284
rect 149900 16282 149906 16284
rect 316217 16282 316283 16285
rect 149900 16280 316283 16282
rect 149900 16224 316222 16280
rect 316278 16224 316283 16280
rect 149900 16222 316283 16224
rect 149900 16220 149906 16222
rect 316217 16219 316283 16222
rect 154246 16084 154252 16148
rect 154316 16146 154322 16148
rect 371233 16146 371299 16149
rect 154316 16144 371299 16146
rect 154316 16088 371238 16144
rect 371294 16088 371299 16144
rect 154316 16086 371299 16088
rect 154316 16084 154322 16086
rect 371233 16083 371299 16086
rect 155718 15948 155724 16012
rect 155788 16010 155794 16012
rect 387793 16010 387859 16013
rect 155788 16008 387859 16010
rect 155788 15952 387798 16008
rect 387854 15952 387859 16008
rect 155788 15950 387859 15952
rect 155788 15948 155794 15950
rect 387793 15947 387859 15950
rect 158294 15812 158300 15876
rect 158364 15874 158370 15876
rect 420913 15874 420979 15877
rect 158364 15872 420979 15874
rect 158364 15816 420918 15872
rect 420974 15816 420979 15872
rect 158364 15814 420979 15816
rect 158364 15812 158370 15814
rect 420913 15811 420979 15814
rect 154430 14724 154436 14788
rect 154500 14786 154506 14788
rect 370129 14786 370195 14789
rect 154500 14784 370195 14786
rect 154500 14728 370134 14784
rect 370190 14728 370195 14784
rect 154500 14726 370195 14728
rect 154500 14724 154506 14726
rect 370129 14723 370195 14726
rect 157006 14588 157012 14652
rect 157076 14650 157082 14652
rect 407205 14650 407271 14653
rect 157076 14648 407271 14650
rect 157076 14592 407210 14648
rect 407266 14592 407271 14648
rect 157076 14590 407271 14592
rect 157076 14588 157082 14590
rect 407205 14587 407271 14590
rect 162526 14452 162532 14516
rect 162596 14514 162602 14516
rect 478137 14514 478203 14517
rect 162596 14512 478203 14514
rect 162596 14456 478142 14512
rect 478198 14456 478203 14512
rect 162596 14454 478203 14456
rect 162596 14452 162602 14454
rect 478137 14451 478203 14454
rect 148542 13228 148548 13292
rect 148612 13290 148618 13292
rect 301497 13290 301563 13293
rect 148612 13288 301563 13290
rect 148612 13232 301502 13288
rect 301558 13232 301563 13288
rect 148612 13230 301563 13232
rect 148612 13228 148618 13230
rect 301497 13227 301563 13230
rect 152958 13092 152964 13156
rect 153028 13154 153034 13156
rect 349245 13154 349311 13157
rect 153028 13152 349311 13154
rect 153028 13096 349250 13152
rect 349306 13096 349311 13152
rect 153028 13094 349311 13096
rect 153028 13092 153034 13094
rect 349245 13091 349311 13094
rect 166758 12956 166764 13020
rect 166828 13018 166834 13020
rect 531405 13018 531471 13021
rect 166828 13016 531471 13018
rect 166828 12960 531410 13016
rect 531466 12960 531471 13016
rect 166828 12958 531471 12960
rect 166828 12956 166834 12958
rect 531405 12955 531471 12958
rect 158478 11732 158484 11796
rect 158548 11794 158554 11796
rect 423765 11794 423831 11797
rect 158548 11792 423831 11794
rect 158548 11736 423770 11792
rect 423826 11736 423831 11792
rect 158548 11734 423831 11736
rect 158548 11732 158554 11734
rect 423765 11731 423831 11734
rect 162710 11596 162716 11660
rect 162780 11658 162786 11660
rect 474089 11658 474155 11661
rect 162780 11656 474155 11658
rect 162780 11600 474094 11656
rect 474150 11600 474155 11656
rect 162780 11598 474155 11600
rect 162780 11596 162786 11598
rect 474089 11595 474155 11598
rect 140998 10644 141004 10708
rect 141068 10706 141074 10708
rect 213361 10706 213427 10709
rect 141068 10704 213427 10706
rect 141068 10648 213366 10704
rect 213422 10648 213427 10704
rect 141068 10646 213427 10648
rect 141068 10644 141074 10646
rect 213361 10643 213427 10646
rect 147070 10508 147076 10572
rect 147140 10570 147146 10572
rect 281533 10570 281599 10573
rect 147140 10568 281599 10570
rect 147140 10512 281538 10568
rect 281594 10512 281599 10568
rect 147140 10510 281599 10512
rect 147140 10508 147146 10510
rect 281533 10507 281599 10510
rect 110505 10434 110571 10437
rect 134190 10434 134196 10436
rect 110505 10432 134196 10434
rect 110505 10376 110510 10432
rect 110566 10376 134196 10432
rect 110505 10374 134196 10376
rect 110505 10371 110571 10374
rect 134190 10372 134196 10374
rect 134260 10372 134266 10436
rect 148726 10372 148732 10436
rect 148796 10434 148802 10436
rect 299657 10434 299723 10437
rect 148796 10432 299723 10434
rect 148796 10376 299662 10432
rect 299718 10376 299723 10432
rect 148796 10374 299723 10376
rect 148796 10372 148802 10374
rect 299657 10371 299723 10374
rect 92473 10298 92539 10301
rect 133086 10298 133092 10300
rect 92473 10296 133092 10298
rect 92473 10240 92478 10296
rect 92534 10240 133092 10296
rect 92473 10238 133092 10240
rect 92473 10235 92539 10238
rect 133086 10236 133092 10238
rect 133156 10236 133162 10300
rect 164918 10236 164924 10300
rect 164988 10298 164994 10300
rect 513373 10298 513439 10301
rect 164988 10296 513439 10298
rect 164988 10240 513378 10296
rect 513434 10240 513439 10296
rect 164988 10238 513439 10240
rect 164988 10236 164994 10238
rect 513373 10235 513439 10238
rect 145414 9148 145420 9212
rect 145484 9210 145490 9212
rect 264145 9210 264211 9213
rect 145484 9208 264211 9210
rect 145484 9152 264150 9208
rect 264206 9152 264211 9208
rect 145484 9150 264211 9152
rect 145484 9148 145490 9150
rect 264145 9147 264211 9150
rect 78581 9074 78647 9077
rect 131430 9074 131436 9076
rect 78581 9072 131436 9074
rect 78581 9016 78586 9072
rect 78642 9016 131436 9072
rect 78581 9014 131436 9016
rect 78581 9011 78647 9014
rect 131430 9012 131436 9014
rect 131500 9012 131506 9076
rect 148358 9012 148364 9076
rect 148428 9074 148434 9076
rect 300761 9074 300827 9077
rect 148428 9072 300827 9074
rect 148428 9016 300766 9072
rect 300822 9016 300827 9072
rect 148428 9014 300827 9016
rect 148428 9012 148434 9014
rect 300761 9011 300827 9014
rect 57145 8938 57211 8941
rect 129958 8938 129964 8940
rect 57145 8936 129964 8938
rect 57145 8880 57150 8936
rect 57206 8880 129964 8936
rect 57145 8878 129964 8880
rect 57145 8875 57211 8878
rect 129958 8876 129964 8878
rect 130028 8876 130034 8940
rect 156638 8876 156644 8940
rect 156708 8938 156714 8940
rect 408401 8938 408467 8941
rect 156708 8936 408467 8938
rect 156708 8880 408406 8936
rect 408462 8880 408467 8936
rect 156708 8878 408467 8880
rect 156708 8876 156714 8878
rect 408401 8875 408467 8878
rect 109309 7986 109375 7989
rect 134006 7986 134012 7988
rect 109309 7984 134012 7986
rect 109309 7928 109314 7984
rect 109370 7928 134012 7984
rect 109309 7926 134012 7928
rect 109309 7923 109375 7926
rect 134006 7924 134012 7926
rect 134076 7924 134082 7988
rect 56041 7850 56107 7853
rect 130142 7850 130148 7852
rect 56041 7848 130148 7850
rect 56041 7792 56046 7848
rect 56102 7792 130148 7848
rect 56041 7790 130148 7792
rect 56041 7787 56107 7790
rect 130142 7788 130148 7790
rect 130212 7788 130218 7852
rect 41873 7714 41939 7717
rect 128670 7714 128676 7716
rect 41873 7712 128676 7714
rect 41873 7656 41878 7712
rect 41934 7656 128676 7712
rect 41873 7654 128676 7656
rect 41873 7651 41939 7654
rect 128670 7652 128676 7654
rect 128740 7652 128746 7716
rect 144310 7652 144316 7716
rect 144380 7714 144386 7716
rect 246389 7714 246455 7717
rect 144380 7712 246455 7714
rect 144380 7656 246394 7712
rect 246450 7656 246455 7712
rect 144380 7654 246455 7656
rect 144380 7652 144386 7654
rect 246389 7651 246455 7654
rect 38377 7578 38443 7581
rect 129038 7578 129044 7580
rect 38377 7576 129044 7578
rect 38377 7520 38382 7576
rect 38438 7520 129044 7576
rect 38377 7518 129044 7520
rect 38377 7515 38443 7518
rect 129038 7516 129044 7518
rect 129108 7516 129114 7580
rect 145598 7516 145604 7580
rect 145668 7578 145674 7580
rect 265341 7578 265407 7581
rect 145668 7576 265407 7578
rect 145668 7520 265346 7576
rect 265402 7520 265407 7576
rect 145668 7518 265407 7520
rect 145668 7516 145674 7518
rect 265341 7515 265407 7518
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 151302 6428 151308 6492
rect 151372 6490 151378 6492
rect 336273 6490 336339 6493
rect 151372 6488 336339 6490
rect 151372 6432 336278 6488
rect 336334 6432 336339 6488
rect 583520 6476 584960 6566
rect 151372 6430 336339 6432
rect 151372 6428 151378 6430
rect 336273 6427 336339 6430
rect 111609 6354 111675 6357
rect 134374 6354 134380 6356
rect 111609 6352 134380 6354
rect 111609 6296 111614 6352
rect 111670 6296 134380 6352
rect 111609 6294 134380 6296
rect 111609 6291 111675 6294
rect 134374 6292 134380 6294
rect 134444 6292 134450 6356
rect 151486 6292 151492 6356
rect 151556 6354 151562 6356
rect 337469 6354 337535 6357
rect 151556 6352 337535 6354
rect 151556 6296 337474 6352
rect 337530 6296 337535 6352
rect 151556 6294 337535 6296
rect 151556 6292 151562 6294
rect 337469 6291 337535 6294
rect 73797 6218 73863 6221
rect 131246 6218 131252 6220
rect 73797 6216 131252 6218
rect 73797 6160 73802 6216
rect 73858 6160 131252 6216
rect 73797 6158 131252 6160
rect 73797 6155 73863 6158
rect 131246 6156 131252 6158
rect 131316 6156 131322 6220
rect 131982 6156 131988 6220
rect 132052 6218 132058 6220
rect 333881 6218 333947 6221
rect 132052 6216 333947 6218
rect 132052 6160 333886 6216
rect 333942 6160 333947 6216
rect 132052 6158 333947 6160
rect 132052 6156 132058 6158
rect 333881 6155 333947 6158
rect 150014 5068 150020 5132
rect 150084 5130 150090 5132
rect 315021 5130 315087 5133
rect 150084 5128 315087 5130
rect 150084 5072 315026 5128
rect 315082 5072 315087 5128
rect 150084 5070 315087 5072
rect 150084 5068 150090 5070
rect 315021 5067 315087 5070
rect 159030 4932 159036 4996
rect 159100 4994 159106 4996
rect 442625 4994 442691 4997
rect 159100 4992 442691 4994
rect 159100 4936 442630 4992
rect 442686 4936 442691 4992
rect 159100 4934 442691 4936
rect 159100 4932 159106 4934
rect 442625 4931 442691 4934
rect 4061 4858 4127 4861
rect 125726 4858 125732 4860
rect 4061 4856 125732 4858
rect 4061 4800 4066 4856
rect 4122 4800 125732 4856
rect 4061 4798 125732 4800
rect 4061 4795 4127 4798
rect 125726 4796 125732 4798
rect 125796 4796 125802 4860
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 158897 4858 158963 4861
rect 137940 4856 158963 4858
rect 137940 4800 158902 4856
rect 158958 4800 158963 4856
rect 137940 4798 158963 4800
rect 137940 4796 137946 4798
rect 158897 4795 158963 4798
rect 168046 4796 168052 4860
rect 168116 4858 168122 4860
rect 547873 4858 547939 4861
rect 168116 4856 547939 4858
rect 168116 4800 547878 4856
rect 547934 4800 547939 4856
rect 168116 4798 547939 4800
rect 168116 4796 168122 4798
rect 547873 4795 547939 4798
rect 151670 3572 151676 3636
rect 151740 3634 151746 3636
rect 335077 3634 335143 3637
rect 151740 3632 335143 3634
rect 151740 3576 335082 3632
rect 335138 3576 335143 3632
rect 151740 3574 335143 3576
rect 151740 3572 151746 3574
rect 335077 3571 335143 3574
rect 72601 3498 72667 3501
rect 131062 3498 131068 3500
rect 72601 3496 131068 3498
rect 72601 3440 72606 3496
rect 72662 3440 131068 3496
rect 72601 3438 131068 3440
rect 72601 3435 72667 3438
rect 131062 3436 131068 3438
rect 131132 3436 131138 3500
rect 171726 3436 171732 3500
rect 171796 3498 171802 3500
rect 570321 3498 570387 3501
rect 171796 3496 570387 3498
rect 171796 3440 570326 3496
rect 570382 3440 570387 3496
rect 171796 3438 570387 3440
rect 171796 3436 171802 3438
rect 570321 3435 570387 3438
rect 20621 3362 20687 3365
rect 127014 3362 127020 3364
rect 20621 3360 127020 3362
rect 20621 3304 20626 3360
rect 20682 3304 127020 3360
rect 20621 3302 127020 3304
rect 20621 3299 20687 3302
rect 127014 3300 127020 3302
rect 127084 3300 127090 3364
rect 136398 3300 136404 3364
rect 136468 3362 136474 3364
rect 161289 3362 161355 3365
rect 136468 3360 161355 3362
rect 136468 3304 161294 3360
rect 161350 3304 161355 3360
rect 136468 3302 161355 3304
rect 136468 3300 136474 3302
rect 161289 3299 161355 3302
rect 171910 3300 171916 3364
rect 171980 3362 171986 3364
rect 580993 3362 581059 3365
rect 171980 3360 581059 3362
rect 171980 3304 580998 3360
rect 581054 3304 581059 3360
rect 171980 3302 581059 3304
rect 171980 3300 171986 3302
rect 580993 3299 581059 3302
<< via3 >>
rect 396580 696900 396644 696964
rect 144500 190980 144564 191044
rect 146156 188532 146220 188596
rect 144500 188124 144564 188188
rect 141188 184316 141252 184380
rect 141004 184180 141068 184244
rect 143028 184044 143092 184108
rect 148732 181188 148796 181252
rect 144684 180976 144748 180980
rect 144684 180920 144698 180976
rect 144698 180920 144748 180976
rect 144684 180916 144748 180920
rect 143028 178876 143092 178940
rect 141188 178740 141252 178804
rect 141004 178604 141068 178668
rect 148732 171804 148796 171868
rect 146156 142836 146220 142900
rect 144684 142700 144748 142764
rect 173388 81228 173452 81292
rect 171180 81092 171244 81156
rect 171916 80956 171980 81020
rect 172100 80684 172164 80748
rect 173020 80548 173084 80612
rect 172836 80412 172900 80476
rect 158668 80140 158732 80204
rect 125732 79928 125796 79932
rect 125732 79872 125736 79928
rect 125736 79872 125792 79928
rect 125792 79872 125796 79928
rect 125732 79868 125796 79872
rect 127020 79868 127084 79932
rect 127204 79732 127268 79796
rect 128676 79906 128680 79932
rect 128680 79906 128736 79932
rect 128736 79906 128740 79932
rect 128676 79868 128740 79906
rect 130332 80004 130396 80068
rect 144684 80004 144748 80068
rect 151492 80004 151556 80068
rect 130516 79868 130580 79932
rect 131252 79906 131256 79932
rect 131256 79906 131312 79932
rect 131312 79906 131316 79932
rect 131252 79868 131316 79906
rect 128860 79732 128924 79796
rect 131620 79906 131624 79932
rect 131624 79906 131680 79932
rect 131680 79906 131684 79932
rect 131620 79868 131684 79906
rect 129044 79596 129108 79660
rect 133276 79868 133340 79932
rect 134196 79906 134200 79932
rect 134200 79906 134256 79932
rect 134256 79906 134260 79932
rect 134196 79868 134260 79906
rect 134012 79792 134076 79796
rect 134012 79736 134016 79792
rect 134016 79736 134072 79792
rect 134072 79736 134076 79792
rect 134012 79732 134076 79736
rect 135300 79732 135364 79796
rect 137692 79868 137756 79932
rect 138428 79906 138432 79932
rect 138432 79906 138488 79932
rect 138488 79906 138492 79932
rect 138428 79868 138492 79906
rect 138612 79732 138676 79796
rect 138980 79732 139044 79796
rect 134196 79596 134260 79660
rect 140452 79868 140516 79932
rect 142476 79868 142540 79932
rect 142844 79868 142908 79932
rect 143028 79732 143092 79796
rect 143764 79868 143828 79932
rect 144132 79732 144196 79796
rect 141004 79596 141068 79660
rect 143212 79656 143276 79660
rect 143212 79600 143262 79656
rect 143262 79600 143276 79656
rect 143212 79596 143276 79600
rect 144500 79732 144564 79796
rect 145972 79928 146036 79932
rect 145972 79872 145976 79928
rect 145976 79872 146032 79928
rect 146032 79872 146036 79928
rect 145972 79868 146036 79872
rect 147260 79868 147324 79932
rect 148180 79868 148244 79932
rect 148916 79868 148980 79932
rect 149100 79868 149164 79932
rect 145604 79732 145668 79796
rect 150388 79894 150452 79932
rect 150388 79868 150392 79894
rect 150392 79868 150448 79894
rect 150448 79868 150452 79894
rect 150756 79868 150820 79932
rect 151308 79906 151312 79932
rect 151312 79906 151368 79932
rect 151368 79906 151372 79932
rect 159772 80140 159836 80204
rect 171364 80276 171428 80340
rect 171548 80276 171612 80340
rect 165108 80140 165172 80204
rect 151308 79868 151372 79906
rect 147444 79732 147508 79796
rect 148364 79732 148428 79796
rect 149468 79596 149532 79660
rect 152780 79732 152844 79796
rect 153148 79732 153212 79796
rect 154252 79868 154316 79932
rect 154620 79868 154684 79932
rect 155356 79868 155420 79932
rect 156460 79868 156524 79932
rect 156828 79868 156892 79932
rect 155540 79596 155604 79660
rect 156644 79732 156708 79796
rect 157932 79868 157996 79932
rect 158484 79732 158548 79796
rect 158852 79732 158916 79796
rect 160324 79868 160388 79932
rect 161060 79868 161124 79932
rect 161796 79868 161860 79932
rect 161980 79928 162044 79932
rect 161980 79872 161984 79928
rect 161984 79872 162040 79928
rect 162040 79872 162044 79928
rect 161980 79868 162044 79872
rect 162348 79868 162412 79932
rect 163452 79868 163516 79932
rect 162532 79596 162596 79660
rect 163268 79596 163332 79660
rect 163452 79596 163516 79660
rect 164556 79906 164560 79932
rect 164560 79906 164616 79932
rect 164616 79906 164620 79932
rect 164556 79868 164620 79906
rect 165292 79906 165296 79932
rect 165296 79906 165352 79932
rect 165352 79906 165356 79932
rect 165292 79868 165356 79906
rect 166948 79868 167012 79932
rect 167316 79928 167380 79932
rect 167316 79872 167320 79928
rect 167320 79872 167376 79928
rect 167376 79872 167380 79928
rect 167316 79868 167380 79872
rect 167684 79928 167748 79932
rect 167684 79872 167688 79928
rect 167688 79872 167744 79928
rect 167744 79872 167748 79928
rect 167684 79868 167748 79872
rect 167868 79928 167932 79932
rect 167868 79872 167872 79928
rect 167872 79872 167928 79928
rect 167928 79872 167932 79928
rect 167868 79868 167932 79872
rect 168420 79928 168484 79932
rect 168420 79872 168424 79928
rect 168424 79872 168480 79928
rect 168480 79872 168484 79928
rect 168420 79868 168484 79872
rect 168788 79906 168792 79932
rect 168792 79906 168848 79932
rect 168848 79906 168852 79932
rect 168788 79868 168852 79906
rect 169156 79868 169220 79932
rect 169524 80004 169588 80068
rect 171732 80140 171796 80204
rect 170812 80004 170876 80068
rect 172836 80004 172900 80068
rect 173020 80004 173084 80068
rect 170076 79906 170080 79932
rect 170080 79906 170136 79932
rect 170136 79906 170140 79932
rect 170076 79868 170140 79906
rect 165660 79732 165724 79796
rect 168052 79732 168116 79796
rect 169892 79732 169956 79796
rect 164188 79656 164252 79660
rect 164188 79600 164238 79656
rect 164238 79600 164252 79656
rect 164188 79596 164252 79600
rect 165844 79596 165908 79660
rect 166764 79596 166828 79660
rect 170444 79656 170508 79660
rect 171180 79928 171244 79932
rect 171180 79872 171184 79928
rect 171184 79872 171240 79928
rect 171240 79872 171244 79928
rect 171180 79868 171244 79872
rect 171916 79868 171980 79932
rect 172284 79928 172348 79932
rect 172284 79872 172288 79928
rect 172288 79872 172344 79928
rect 172344 79872 172348 79928
rect 172284 79868 172348 79872
rect 172468 79928 172532 79932
rect 172468 79872 172472 79928
rect 172472 79872 172528 79928
rect 172528 79872 172532 79928
rect 172468 79868 172532 79872
rect 170996 79732 171060 79796
rect 172100 79732 172164 79796
rect 172468 79732 172532 79796
rect 170444 79600 170494 79656
rect 170494 79600 170508 79656
rect 170444 79596 170508 79600
rect 173388 79052 173452 79116
rect 173204 78916 173268 78980
rect 138428 78780 138492 78844
rect 145972 78840 146036 78844
rect 145972 78784 145986 78840
rect 145986 78784 146036 78840
rect 145972 78780 146036 78784
rect 148548 78780 148612 78844
rect 150388 78780 150452 78844
rect 151308 78840 151372 78844
rect 151308 78784 151358 78840
rect 151358 78784 151372 78840
rect 151308 78780 151372 78784
rect 165476 78840 165540 78844
rect 165476 78784 165490 78840
rect 165490 78784 165540 78840
rect 165476 78780 165540 78784
rect 168420 78780 168484 78844
rect 172100 78780 172164 78844
rect 144316 78644 144380 78708
rect 145236 78644 145300 78708
rect 147076 78644 147140 78708
rect 148732 78704 148796 78708
rect 148732 78648 148782 78704
rect 148782 78648 148796 78704
rect 148732 78644 148796 78648
rect 149100 78704 149164 78708
rect 149100 78648 149114 78704
rect 149114 78648 149164 78704
rect 149100 78644 149164 78648
rect 149652 78644 149716 78708
rect 150756 78644 150820 78708
rect 151676 78644 151740 78708
rect 153884 78644 153948 78708
rect 159036 78644 159100 78708
rect 160324 78704 160388 78708
rect 160324 78648 160338 78704
rect 160338 78648 160388 78704
rect 160324 78644 160388 78648
rect 161244 78644 161308 78708
rect 161796 78644 161860 78708
rect 162164 78644 162228 78708
rect 162716 78704 162780 78708
rect 162716 78648 162730 78704
rect 162730 78648 162780 78704
rect 162716 78644 162780 78648
rect 165660 78704 165724 78708
rect 165660 78648 165674 78704
rect 165674 78648 165724 78704
rect 165660 78644 165724 78648
rect 165844 78704 165908 78708
rect 165844 78648 165858 78704
rect 165858 78648 165908 78704
rect 165844 78644 165908 78648
rect 166396 78644 166460 78708
rect 167684 78644 167748 78708
rect 170076 78644 170140 78708
rect 170444 78644 170508 78708
rect 171548 78644 171612 78708
rect 145420 78508 145484 78572
rect 149836 78508 149900 78572
rect 151308 78508 151372 78572
rect 158668 78508 158732 78572
rect 161060 78508 161124 78572
rect 164924 78508 164988 78572
rect 167868 78508 167932 78572
rect 169524 78568 169588 78572
rect 169524 78512 169574 78568
rect 169574 78512 169588 78568
rect 169524 78508 169588 78512
rect 170996 78508 171060 78572
rect 150020 78372 150084 78436
rect 160876 78372 160940 78436
rect 396580 78372 396644 78436
rect 128676 78100 128740 78164
rect 129964 78160 130028 78164
rect 129964 78104 130014 78160
rect 130014 78104 130028 78160
rect 129964 78100 130028 78104
rect 137876 78160 137940 78164
rect 137876 78104 137890 78160
rect 137890 78104 137940 78160
rect 137876 78100 137940 78104
rect 155356 78100 155420 78164
rect 158300 78100 158364 78164
rect 159772 78100 159836 78164
rect 167316 78100 167380 78164
rect 167684 78100 167748 78164
rect 168788 78100 168852 78164
rect 169156 78100 169220 78164
rect 169524 78100 169588 78164
rect 128676 78024 128740 78028
rect 128676 77968 128726 78024
rect 128726 77968 128740 78024
rect 128676 77964 128740 77968
rect 129780 78024 129844 78028
rect 129780 77968 129794 78024
rect 129794 77968 129844 78024
rect 129780 77964 129844 77968
rect 130148 78024 130212 78028
rect 130148 77968 130162 78024
rect 130162 77968 130212 78024
rect 130148 77964 130212 77968
rect 130516 78024 130580 78028
rect 130516 77968 130530 78024
rect 130530 77968 130580 78024
rect 130516 77964 130580 77968
rect 131068 78024 131132 78028
rect 131068 77968 131082 78024
rect 131082 77968 131132 78024
rect 131068 77964 131132 77968
rect 135668 77964 135732 78028
rect 136404 77964 136468 78028
rect 158116 77964 158180 78028
rect 171364 77828 171428 77892
rect 131988 77556 132052 77620
rect 163084 77692 163148 77756
rect 163268 77556 163332 77620
rect 164556 77556 164620 77620
rect 166764 77616 166828 77620
rect 166764 77560 166814 77616
rect 166814 77560 166828 77616
rect 166764 77556 166828 77560
rect 168052 77616 168116 77620
rect 168052 77560 168102 77616
rect 168102 77560 168116 77616
rect 168052 77556 168116 77560
rect 133092 77420 133156 77484
rect 148180 77420 148244 77484
rect 157012 77480 157076 77484
rect 157012 77424 157062 77480
rect 157062 77424 157076 77480
rect 157012 77420 157076 77424
rect 152596 77284 152660 77348
rect 161980 77148 162044 77212
rect 172284 77284 172348 77348
rect 172468 77148 172532 77212
rect 142476 77012 142540 77076
rect 152964 76604 153028 76668
rect 128860 76468 128924 76532
rect 169892 76332 169956 76396
rect 155724 76196 155788 76260
rect 142844 76060 142908 76124
rect 125732 75984 125796 75988
rect 125732 75928 125782 75984
rect 125782 75928 125796 75984
rect 125732 75924 125796 75928
rect 140268 75924 140332 75988
rect 142844 75924 142908 75988
rect 143764 75984 143828 75988
rect 143764 75928 143814 75984
rect 143814 75928 143828 75984
rect 143764 75924 143828 75928
rect 154436 75984 154500 75988
rect 154436 75928 154450 75984
rect 154450 75928 154500 75984
rect 154436 75924 154500 75928
rect 154620 75924 154684 75988
rect 156460 75924 156524 75988
rect 171916 75924 171980 75988
rect 140084 75788 140148 75852
rect 154068 75788 154132 75852
rect 130332 75516 130396 75580
rect 129780 75380 129844 75444
rect 125548 75108 125612 75172
rect 167132 75108 167196 75172
rect 135300 74428 135364 74492
rect 144132 73884 144196 73948
rect 144684 73748 144748 73812
rect 162164 72660 162228 72724
rect 147444 72524 147508 72588
rect 148916 72388 148980 72452
rect 153148 71164 153212 71228
rect 163452 71028 163516 71092
rect 138980 69532 139044 69596
rect 165476 68172 165540 68236
rect 140268 65452 140332 65516
rect 166396 62868 166460 62932
rect 172100 62732 172164 62796
rect 160692 61372 160756 61436
rect 138612 60012 138676 60076
rect 143028 59876 143092 59940
rect 149468 53076 149532 53140
rect 152596 47500 152660 47564
rect 135668 44916 135732 44980
rect 133276 44780 133340 44844
rect 147260 44780 147324 44844
rect 127204 43420 127268 43484
rect 153884 40564 153948 40628
rect 154068 35124 154132 35188
rect 143212 34036 143276 34100
rect 145236 33900 145300 33964
rect 170628 33764 170692 33828
rect 166580 32540 166644 32604
rect 169524 32404 169588 32468
rect 167684 30908 167748 30972
rect 149652 29548 149716 29612
rect 140452 28460 140516 28524
rect 142844 28324 142908 28388
rect 165108 28188 165172 28252
rect 165292 26964 165356 27028
rect 170812 26828 170876 26892
rect 155540 25468 155604 25532
rect 157932 24108 157996 24172
rect 170444 21660 170508 21724
rect 158852 21524 158916 21588
rect 160876 21388 160940 21452
rect 162348 21252 162412 21316
rect 144500 20164 144564 20228
rect 161060 20028 161124 20092
rect 137692 19892 137756 19956
rect 163636 19892 163700 19956
rect 140084 18940 140148 19004
rect 152780 18804 152844 18868
rect 158116 18668 158180 18732
rect 167868 18532 167932 18596
rect 156828 17308 156892 17372
rect 161244 17172 161308 17236
rect 149836 16220 149900 16284
rect 154252 16084 154316 16148
rect 155724 15948 155788 16012
rect 158300 15812 158364 15876
rect 154436 14724 154500 14788
rect 157012 14588 157076 14652
rect 162532 14452 162596 14516
rect 148548 13228 148612 13292
rect 152964 13092 153028 13156
rect 166764 12956 166828 13020
rect 158484 11732 158548 11796
rect 162716 11596 162780 11660
rect 141004 10644 141068 10708
rect 147076 10508 147140 10572
rect 134196 10372 134260 10436
rect 148732 10372 148796 10436
rect 133092 10236 133156 10300
rect 164924 10236 164988 10300
rect 145420 9148 145484 9212
rect 131436 9012 131500 9076
rect 148364 9012 148428 9076
rect 129964 8876 130028 8940
rect 156644 8876 156708 8940
rect 134012 7924 134076 7988
rect 130148 7788 130212 7852
rect 128676 7652 128740 7716
rect 144316 7652 144380 7716
rect 129044 7516 129108 7580
rect 145604 7516 145668 7580
rect 151308 6428 151372 6492
rect 134380 6292 134444 6356
rect 151492 6292 151556 6356
rect 131252 6156 131316 6220
rect 131988 6156 132052 6220
rect 150020 5068 150084 5132
rect 159036 4932 159100 4996
rect 125732 4796 125796 4860
rect 137876 4796 137940 4860
rect 168052 4796 168116 4860
rect 151676 3572 151740 3636
rect 131068 3436 131132 3500
rect 171732 3436 171796 3500
rect 127020 3300 127084 3364
rect 136404 3300 136468 3364
rect 171916 3300 171980 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 396579 696964 396645 696965
rect 396579 696900 396580 696964
rect 396644 696900 396645 696964
rect 396579 696899 396645 696900
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 144499 191044 144565 191045
rect 144499 190980 144500 191044
rect 144564 190980 144565 191044
rect 144499 190979 144565 190980
rect 144502 188189 144562 190979
rect 146155 188596 146221 188597
rect 146155 188532 146156 188596
rect 146220 188532 146221 188596
rect 146155 188531 146221 188532
rect 144499 188188 144565 188189
rect 144499 188124 144500 188188
rect 144564 188124 144565 188188
rect 144499 188123 144565 188124
rect 141187 184380 141253 184381
rect 141187 184316 141188 184380
rect 141252 184316 141253 184380
rect 141187 184315 141253 184316
rect 141003 184244 141069 184245
rect 141003 184180 141004 184244
rect 141068 184180 141069 184244
rect 141003 184179 141069 184180
rect 141006 178669 141066 184179
rect 141190 178805 141250 184315
rect 143027 184108 143093 184109
rect 143027 184044 143028 184108
rect 143092 184044 143093 184108
rect 143027 184043 143093 184044
rect 143030 178941 143090 184043
rect 144683 180980 144749 180981
rect 144683 180916 144684 180980
rect 144748 180916 144749 180980
rect 144683 180915 144749 180916
rect 143027 178940 143093 178941
rect 143027 178876 143028 178940
rect 143092 178876 143093 178940
rect 143027 178875 143093 178876
rect 141187 178804 141253 178805
rect 141187 178740 141188 178804
rect 141252 178740 141253 178804
rect 141187 178739 141253 178740
rect 141003 178668 141069 178669
rect 141003 178604 141004 178668
rect 141068 178604 141069 178668
rect 141003 178603 141069 178604
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 144686 142765 144746 180915
rect 146158 142901 146218 188531
rect 148731 181252 148797 181253
rect 148731 181188 148732 181252
rect 148796 181188 148797 181252
rect 148731 181187 148797 181188
rect 148734 171869 148794 181187
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 148731 171868 148797 171869
rect 148731 171804 148732 171868
rect 148796 171804 148797 171868
rect 148731 171803 148797 171804
rect 146155 142900 146221 142901
rect 146155 142836 146156 142900
rect 146220 142836 146221 142900
rect 146155 142835 146221 142836
rect 144683 142764 144749 142765
rect 144683 142700 144684 142764
rect 144748 142700 144749 142764
rect 144683 142699 144749 142700
rect 172794 142000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 173387 81292 173453 81293
rect 173387 81228 173388 81292
rect 173452 81228 173453 81292
rect 173387 81227 173453 81228
rect 171179 81156 171245 81157
rect 171179 81092 171180 81156
rect 171244 81092 171245 81156
rect 171179 81091 171245 81092
rect 158667 80204 158733 80205
rect 158667 80140 158668 80204
rect 158732 80140 158733 80204
rect 158667 80139 158733 80140
rect 159771 80204 159837 80205
rect 159771 80140 159772 80204
rect 159836 80140 159837 80204
rect 159771 80139 159837 80140
rect 165107 80204 165173 80205
rect 165107 80140 165108 80204
rect 165172 80140 165173 80204
rect 165107 80139 165173 80140
rect 130331 80068 130397 80069
rect 130331 80004 130332 80068
rect 130396 80004 130397 80068
rect 130331 80003 130397 80004
rect 144683 80068 144749 80069
rect 144683 80004 144684 80068
rect 144748 80004 144749 80068
rect 144683 80003 144749 80004
rect 151491 80068 151557 80069
rect 151491 80004 151492 80068
rect 151556 80004 151557 80068
rect 151491 80003 151557 80004
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 125731 79932 125797 79933
rect 125731 79930 125732 79932
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 125550 79870 125732 79930
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125550 75173 125610 79870
rect 125731 79868 125732 79870
rect 125796 79868 125797 79932
rect 125731 79867 125797 79868
rect 127019 79932 127085 79933
rect 127019 79868 127020 79932
rect 127084 79868 127085 79932
rect 127019 79867 127085 79868
rect 128675 79932 128741 79933
rect 128675 79868 128676 79932
rect 128740 79868 128741 79932
rect 128675 79867 128741 79868
rect 125731 75988 125797 75989
rect 125731 75924 125732 75988
rect 125796 75924 125797 75988
rect 125731 75923 125797 75924
rect 125547 75172 125613 75173
rect 125547 75108 125548 75172
rect 125612 75108 125613 75172
rect 125547 75107 125613 75108
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 125734 4861 125794 75923
rect 125731 4860 125797 4861
rect 125731 4796 125732 4860
rect 125796 4796 125797 4860
rect 125731 4795 125797 4796
rect 127022 3365 127082 79867
rect 127203 79796 127269 79797
rect 127203 79732 127204 79796
rect 127268 79732 127269 79796
rect 127203 79731 127269 79732
rect 127206 43485 127266 79731
rect 128678 78165 128738 79867
rect 128859 79796 128925 79797
rect 128859 79732 128860 79796
rect 128924 79732 128925 79796
rect 128859 79731 128925 79732
rect 128675 78164 128741 78165
rect 128675 78100 128676 78164
rect 128740 78100 128741 78164
rect 128675 78099 128741 78100
rect 128675 78028 128741 78029
rect 127794 57454 128414 78000
rect 128675 77964 128676 78028
rect 128740 77964 128741 78028
rect 128675 77963 128741 77964
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127203 43484 127269 43485
rect 127203 43420 127204 43484
rect 127268 43420 127269 43484
rect 127203 43419 127269 43420
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127019 3364 127085 3365
rect 127019 3300 127020 3364
rect 127084 3300 127085 3364
rect 127019 3299 127085 3300
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128678 7717 128738 77963
rect 128862 76533 128922 79731
rect 129043 79660 129109 79661
rect 129043 79596 129044 79660
rect 129108 79596 129109 79660
rect 129043 79595 129109 79596
rect 128859 76532 128925 76533
rect 128859 76468 128860 76532
rect 128924 76468 128925 76532
rect 128859 76467 128925 76468
rect 128675 7716 128741 7717
rect 128675 7652 128676 7716
rect 128740 7652 128741 7716
rect 128675 7651 128741 7652
rect 129046 7581 129106 79595
rect 129963 78164 130029 78165
rect 129963 78100 129964 78164
rect 130028 78100 130029 78164
rect 129963 78099 130029 78100
rect 129779 78028 129845 78029
rect 129779 77964 129780 78028
rect 129844 77964 129845 78028
rect 129779 77963 129845 77964
rect 129782 75445 129842 77963
rect 129779 75444 129845 75445
rect 129779 75380 129780 75444
rect 129844 75380 129845 75444
rect 129779 75379 129845 75380
rect 129966 8941 130026 78099
rect 130147 78028 130213 78029
rect 130147 77964 130148 78028
rect 130212 77964 130213 78028
rect 130147 77963 130213 77964
rect 129963 8940 130029 8941
rect 129963 8876 129964 8940
rect 130028 8876 130029 8940
rect 129963 8875 130029 8876
rect 130150 7853 130210 77963
rect 130334 75581 130394 80003
rect 130515 79932 130581 79933
rect 130515 79868 130516 79932
rect 130580 79868 130581 79932
rect 130515 79867 130581 79868
rect 131251 79932 131317 79933
rect 131251 79868 131252 79932
rect 131316 79868 131317 79932
rect 131251 79867 131317 79868
rect 131619 79932 131685 79933
rect 131619 79868 131620 79932
rect 131684 79868 131685 79932
rect 131619 79867 131685 79868
rect 133275 79932 133341 79933
rect 133275 79868 133276 79932
rect 133340 79868 133341 79932
rect 133275 79867 133341 79868
rect 134195 79932 134261 79933
rect 134195 79868 134196 79932
rect 134260 79930 134261 79932
rect 137691 79932 137757 79933
rect 134260 79870 134442 79930
rect 134260 79868 134261 79870
rect 134195 79867 134261 79868
rect 130518 78029 130578 79867
rect 130515 78028 130581 78029
rect 130515 77964 130516 78028
rect 130580 77964 130581 78028
rect 130515 77963 130581 77964
rect 131067 78028 131133 78029
rect 131067 77964 131068 78028
rect 131132 77964 131133 78028
rect 131067 77963 131133 77964
rect 130331 75580 130397 75581
rect 130331 75516 130332 75580
rect 130396 75516 130397 75580
rect 130331 75515 130397 75516
rect 130147 7852 130213 7853
rect 130147 7788 130148 7852
rect 130212 7788 130213 7852
rect 130147 7787 130213 7788
rect 129043 7580 129109 7581
rect 129043 7516 129044 7580
rect 129108 7516 129109 7580
rect 129043 7515 129109 7516
rect 131070 3501 131130 77963
rect 131254 6221 131314 79867
rect 131622 75930 131682 79867
rect 131987 77620 132053 77621
rect 131987 77556 131988 77620
rect 132052 77556 132053 77620
rect 131987 77555 132053 77556
rect 131438 75870 131682 75930
rect 131438 9077 131498 75870
rect 131435 9076 131501 9077
rect 131435 9012 131436 9076
rect 131500 9012 131501 9076
rect 131435 9011 131501 9012
rect 131990 6221 132050 77555
rect 132294 61954 132914 78000
rect 133091 77484 133157 77485
rect 133091 77420 133092 77484
rect 133156 77420 133157 77484
rect 133091 77419 133157 77420
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131251 6220 131317 6221
rect 131251 6156 131252 6220
rect 131316 6156 131317 6220
rect 131251 6155 131317 6156
rect 131987 6220 132053 6221
rect 131987 6156 131988 6220
rect 132052 6156 132053 6220
rect 131987 6155 132053 6156
rect 131067 3500 131133 3501
rect 131067 3436 131068 3500
rect 131132 3436 131133 3500
rect 131067 3435 131133 3436
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 10301 133154 77419
rect 133278 44845 133338 79867
rect 134011 79796 134077 79797
rect 134011 79732 134012 79796
rect 134076 79732 134077 79796
rect 134011 79731 134077 79732
rect 133275 44844 133341 44845
rect 133275 44780 133276 44844
rect 133340 44780 133341 44844
rect 133275 44779 133341 44780
rect 133091 10300 133157 10301
rect 133091 10236 133092 10300
rect 133156 10236 133157 10300
rect 133091 10235 133157 10236
rect 134014 7989 134074 79731
rect 134195 79660 134261 79661
rect 134195 79596 134196 79660
rect 134260 79596 134261 79660
rect 134195 79595 134261 79596
rect 134198 10437 134258 79595
rect 134195 10436 134261 10437
rect 134195 10372 134196 10436
rect 134260 10372 134261 10436
rect 134195 10371 134261 10372
rect 134011 7988 134077 7989
rect 134011 7924 134012 7988
rect 134076 7924 134077 7988
rect 134011 7923 134077 7924
rect 134382 6357 134442 79870
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138427 79932 138493 79933
rect 138427 79868 138428 79932
rect 138492 79868 138493 79932
rect 138427 79867 138493 79868
rect 140451 79932 140517 79933
rect 140451 79868 140452 79932
rect 140516 79868 140517 79932
rect 140451 79867 140517 79868
rect 142475 79932 142541 79933
rect 142475 79868 142476 79932
rect 142540 79868 142541 79932
rect 142475 79867 142541 79868
rect 142843 79932 142909 79933
rect 142843 79868 142844 79932
rect 142908 79868 142909 79932
rect 142843 79867 142909 79868
rect 143763 79932 143829 79933
rect 143763 79868 143764 79932
rect 143828 79868 143829 79932
rect 143763 79867 143829 79868
rect 135299 79796 135365 79797
rect 135299 79732 135300 79796
rect 135364 79732 135365 79796
rect 135299 79731 135365 79732
rect 135302 74493 135362 79731
rect 135667 78028 135733 78029
rect 135667 77964 135668 78028
rect 135732 77964 135733 78028
rect 135667 77963 135733 77964
rect 136403 78028 136469 78029
rect 136403 77964 136404 78028
rect 136468 77964 136469 78028
rect 136403 77963 136469 77964
rect 135299 74492 135365 74493
rect 135299 74428 135300 74492
rect 135364 74428 135365 74492
rect 135299 74427 135365 74428
rect 135670 44981 135730 77963
rect 135667 44980 135733 44981
rect 135667 44916 135668 44980
rect 135732 44916 135733 44980
rect 135667 44915 135733 44916
rect 134379 6356 134445 6357
rect 134379 6292 134380 6356
rect 134444 6292 134445 6356
rect 134379 6291 134445 6292
rect 136406 3365 136466 77963
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 3364 136469 3365
rect 136403 3300 136404 3364
rect 136468 3300 136469 3364
rect 136403 3299 136469 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137694 19957 137754 79867
rect 138430 78845 138490 79867
rect 138611 79796 138677 79797
rect 138611 79732 138612 79796
rect 138676 79732 138677 79796
rect 138611 79731 138677 79732
rect 138979 79796 139045 79797
rect 138979 79732 138980 79796
rect 139044 79732 139045 79796
rect 138979 79731 139045 79732
rect 138427 78844 138493 78845
rect 138427 78780 138428 78844
rect 138492 78780 138493 78844
rect 138427 78779 138493 78780
rect 137875 78164 137941 78165
rect 137875 78100 137876 78164
rect 137940 78100 137941 78164
rect 137875 78099 137941 78100
rect 137691 19956 137757 19957
rect 137691 19892 137692 19956
rect 137756 19892 137757 19956
rect 137691 19891 137757 19892
rect 137878 4861 137938 78099
rect 138614 60077 138674 79731
rect 138982 69597 139042 79731
rect 140267 75988 140333 75989
rect 140267 75924 140268 75988
rect 140332 75924 140333 75988
rect 140267 75923 140333 75924
rect 140083 75852 140149 75853
rect 140083 75788 140084 75852
rect 140148 75788 140149 75852
rect 140083 75787 140149 75788
rect 138979 69596 139045 69597
rect 138979 69532 138980 69596
rect 139044 69532 139045 69596
rect 138979 69531 139045 69532
rect 138611 60076 138677 60077
rect 138611 60012 138612 60076
rect 138676 60012 138677 60076
rect 138611 60011 138677 60012
rect 140086 19005 140146 75787
rect 140270 65517 140330 75923
rect 140267 65516 140333 65517
rect 140267 65452 140268 65516
rect 140332 65452 140333 65516
rect 140267 65451 140333 65452
rect 140454 28525 140514 79867
rect 141003 79660 141069 79661
rect 141003 79596 141004 79660
rect 141068 79596 141069 79660
rect 141003 79595 141069 79596
rect 140451 28524 140517 28525
rect 140451 28460 140452 28524
rect 140516 28460 140517 28524
rect 140451 28459 140517 28460
rect 140083 19004 140149 19005
rect 140083 18940 140084 19004
rect 140148 18940 140149 19004
rect 140083 18939 140149 18940
rect 141006 10709 141066 79595
rect 141294 70954 141914 78000
rect 142478 77077 142538 79867
rect 142475 77076 142541 77077
rect 142475 77012 142476 77076
rect 142540 77012 142541 77076
rect 142475 77011 142541 77012
rect 142846 76125 142906 79867
rect 143027 79796 143093 79797
rect 143027 79732 143028 79796
rect 143092 79732 143093 79796
rect 143027 79731 143093 79732
rect 142843 76124 142909 76125
rect 142843 76060 142844 76124
rect 142908 76060 142909 76124
rect 142843 76059 142909 76060
rect 142843 75988 142909 75989
rect 142843 75924 142844 75988
rect 142908 75924 142909 75988
rect 142843 75923 142909 75924
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 10708 141069 10709
rect 141003 10644 141004 10708
rect 141068 10644 141069 10708
rect 141003 10643 141069 10644
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 28389 142906 75923
rect 143030 59941 143090 79731
rect 143211 79660 143277 79661
rect 143211 79596 143212 79660
rect 143276 79596 143277 79660
rect 143211 79595 143277 79596
rect 143027 59940 143093 59941
rect 143027 59876 143028 59940
rect 143092 59876 143093 59940
rect 143027 59875 143093 59876
rect 143214 34101 143274 79595
rect 143766 75989 143826 79867
rect 144131 79796 144197 79797
rect 144131 79732 144132 79796
rect 144196 79732 144197 79796
rect 144131 79731 144197 79732
rect 144499 79796 144565 79797
rect 144499 79732 144500 79796
rect 144564 79732 144565 79796
rect 144499 79731 144565 79732
rect 143763 75988 143829 75989
rect 143763 75924 143764 75988
rect 143828 75924 143829 75988
rect 143763 75923 143829 75924
rect 144134 73949 144194 79731
rect 144315 78708 144381 78709
rect 144315 78644 144316 78708
rect 144380 78644 144381 78708
rect 144315 78643 144381 78644
rect 144131 73948 144197 73949
rect 144131 73884 144132 73948
rect 144196 73884 144197 73948
rect 144131 73883 144197 73884
rect 143211 34100 143277 34101
rect 143211 34036 143212 34100
rect 143276 34036 143277 34100
rect 143211 34035 143277 34036
rect 142843 28388 142909 28389
rect 142843 28324 142844 28388
rect 142908 28324 142909 28388
rect 142843 28323 142909 28324
rect 144318 7717 144378 78643
rect 144502 20229 144562 79731
rect 144686 73813 144746 80003
rect 145971 79932 146037 79933
rect 145971 79868 145972 79932
rect 146036 79868 146037 79932
rect 145971 79867 146037 79868
rect 147259 79932 147325 79933
rect 147259 79868 147260 79932
rect 147324 79868 147325 79932
rect 147259 79867 147325 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148179 79867 148245 79868
rect 148915 79932 148981 79933
rect 148915 79868 148916 79932
rect 148980 79868 148981 79932
rect 148915 79867 148981 79868
rect 149099 79932 149165 79933
rect 149099 79868 149100 79932
rect 149164 79868 149165 79932
rect 149099 79867 149165 79868
rect 150387 79932 150453 79933
rect 150387 79868 150388 79932
rect 150452 79868 150453 79932
rect 150387 79867 150453 79868
rect 150755 79932 150821 79933
rect 150755 79868 150756 79932
rect 150820 79868 150821 79932
rect 150755 79867 150821 79868
rect 151307 79932 151373 79933
rect 151307 79868 151308 79932
rect 151372 79868 151373 79932
rect 151307 79867 151373 79868
rect 145603 79796 145669 79797
rect 145603 79732 145604 79796
rect 145668 79732 145669 79796
rect 145603 79731 145669 79732
rect 145235 78708 145301 78709
rect 145235 78644 145236 78708
rect 145300 78644 145301 78708
rect 145235 78643 145301 78644
rect 144683 73812 144749 73813
rect 144683 73748 144684 73812
rect 144748 73748 144749 73812
rect 144683 73747 144749 73748
rect 145238 33965 145298 78643
rect 145419 78572 145485 78573
rect 145419 78508 145420 78572
rect 145484 78508 145485 78572
rect 145419 78507 145485 78508
rect 145235 33964 145301 33965
rect 145235 33900 145236 33964
rect 145300 33900 145301 33964
rect 145235 33899 145301 33900
rect 144499 20228 144565 20229
rect 144499 20164 144500 20228
rect 144564 20164 144565 20228
rect 144499 20163 144565 20164
rect 145422 9213 145482 78507
rect 145419 9212 145485 9213
rect 145419 9148 145420 9212
rect 145484 9148 145485 9212
rect 145419 9147 145485 9148
rect 144315 7716 144381 7717
rect 144315 7652 144316 7716
rect 144380 7652 144381 7716
rect 144315 7651 144381 7652
rect 145606 7581 145666 79731
rect 145974 78845 146034 79867
rect 145971 78844 146037 78845
rect 145971 78780 145972 78844
rect 146036 78780 146037 78844
rect 145971 78779 146037 78780
rect 147075 78708 147141 78709
rect 147075 78644 147076 78708
rect 147140 78644 147141 78708
rect 147075 78643 147141 78644
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 7580 145669 7581
rect 145603 7516 145604 7580
rect 145668 7516 145669 7580
rect 145603 7515 145669 7516
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 147078 10573 147138 78643
rect 147262 44845 147322 79867
rect 147443 79796 147509 79797
rect 147443 79732 147444 79796
rect 147508 79732 147509 79796
rect 147443 79731 147509 79732
rect 147446 72589 147506 79731
rect 148182 77485 148242 79867
rect 148363 79796 148429 79797
rect 148363 79732 148364 79796
rect 148428 79732 148429 79796
rect 148363 79731 148429 79732
rect 148179 77484 148245 77485
rect 148179 77420 148180 77484
rect 148244 77420 148245 77484
rect 148179 77419 148245 77420
rect 147443 72588 147509 72589
rect 147443 72524 147444 72588
rect 147508 72524 147509 72588
rect 147443 72523 147509 72524
rect 147259 44844 147325 44845
rect 147259 44780 147260 44844
rect 147324 44780 147325 44844
rect 147259 44779 147325 44780
rect 147075 10572 147141 10573
rect 147075 10508 147076 10572
rect 147140 10508 147141 10572
rect 147075 10507 147141 10508
rect 148366 9077 148426 79731
rect 148547 78844 148613 78845
rect 148547 78780 148548 78844
rect 148612 78780 148613 78844
rect 148547 78779 148613 78780
rect 148550 13293 148610 78779
rect 148731 78708 148797 78709
rect 148731 78644 148732 78708
rect 148796 78644 148797 78708
rect 148731 78643 148797 78644
rect 148547 13292 148613 13293
rect 148547 13228 148548 13292
rect 148612 13228 148613 13292
rect 148547 13227 148613 13228
rect 148734 10437 148794 78643
rect 148918 72453 148978 79867
rect 149102 78709 149162 79867
rect 149467 79660 149533 79661
rect 149467 79596 149468 79660
rect 149532 79596 149533 79660
rect 149467 79595 149533 79596
rect 149099 78708 149165 78709
rect 149099 78644 149100 78708
rect 149164 78644 149165 78708
rect 149099 78643 149165 78644
rect 148915 72452 148981 72453
rect 148915 72388 148916 72452
rect 148980 72388 148981 72452
rect 148915 72387 148981 72388
rect 149470 53141 149530 79595
rect 150390 78845 150450 79867
rect 150387 78844 150453 78845
rect 150387 78780 150388 78844
rect 150452 78780 150453 78844
rect 150387 78779 150453 78780
rect 150758 78709 150818 79867
rect 151310 78845 151370 79867
rect 151307 78844 151373 78845
rect 151307 78780 151308 78844
rect 151372 78780 151373 78844
rect 151307 78779 151373 78780
rect 149651 78708 149717 78709
rect 149651 78644 149652 78708
rect 149716 78644 149717 78708
rect 149651 78643 149717 78644
rect 150755 78708 150821 78709
rect 150755 78644 150756 78708
rect 150820 78644 150821 78708
rect 150755 78643 150821 78644
rect 149467 53140 149533 53141
rect 149467 53076 149468 53140
rect 149532 53076 149533 53140
rect 149467 53075 149533 53076
rect 149654 29613 149714 78643
rect 149835 78572 149901 78573
rect 149835 78508 149836 78572
rect 149900 78508 149901 78572
rect 149835 78507 149901 78508
rect 151307 78572 151373 78573
rect 151307 78508 151308 78572
rect 151372 78508 151373 78572
rect 151307 78507 151373 78508
rect 149651 29612 149717 29613
rect 149651 29548 149652 29612
rect 149716 29548 149717 29612
rect 149651 29547 149717 29548
rect 149838 16285 149898 78507
rect 150019 78436 150085 78437
rect 150019 78372 150020 78436
rect 150084 78372 150085 78436
rect 150019 78371 150085 78372
rect 149835 16284 149901 16285
rect 149835 16220 149836 16284
rect 149900 16220 149901 16284
rect 149835 16219 149901 16220
rect 148731 10436 148797 10437
rect 148731 10372 148732 10436
rect 148796 10372 148797 10436
rect 148731 10371 148797 10372
rect 148363 9076 148429 9077
rect 148363 9012 148364 9076
rect 148428 9012 148429 9076
rect 148363 9011 148429 9012
rect 150022 5133 150082 78371
rect 150294 43954 150914 78000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150019 5132 150085 5133
rect 150019 5068 150020 5132
rect 150084 5068 150085 5132
rect 150019 5067 150085 5068
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 151310 6493 151370 78507
rect 151307 6492 151373 6493
rect 151307 6428 151308 6492
rect 151372 6428 151373 6492
rect 151307 6427 151373 6428
rect 151494 6357 151554 80003
rect 154251 79932 154317 79933
rect 154251 79868 154252 79932
rect 154316 79868 154317 79932
rect 154251 79867 154317 79868
rect 154619 79932 154685 79933
rect 154619 79868 154620 79932
rect 154684 79868 154685 79932
rect 154619 79867 154685 79868
rect 155355 79932 155421 79933
rect 155355 79868 155356 79932
rect 155420 79868 155421 79932
rect 155355 79867 155421 79868
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 156459 79867 156525 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79868 156893 79932
rect 156827 79867 156893 79868
rect 157931 79932 157997 79933
rect 157931 79868 157932 79932
rect 157996 79868 157997 79932
rect 157931 79867 157997 79868
rect 152779 79796 152845 79797
rect 152779 79732 152780 79796
rect 152844 79732 152845 79796
rect 152779 79731 152845 79732
rect 153147 79796 153213 79797
rect 153147 79732 153148 79796
rect 153212 79732 153213 79796
rect 153147 79731 153213 79732
rect 151675 78708 151741 78709
rect 151675 78644 151676 78708
rect 151740 78644 151741 78708
rect 151675 78643 151741 78644
rect 151491 6356 151557 6357
rect 151491 6292 151492 6356
rect 151556 6292 151557 6356
rect 151491 6291 151557 6292
rect 151678 3637 151738 78643
rect 152595 77348 152661 77349
rect 152595 77284 152596 77348
rect 152660 77284 152661 77348
rect 152595 77283 152661 77284
rect 152598 47565 152658 77283
rect 152595 47564 152661 47565
rect 152595 47500 152596 47564
rect 152660 47500 152661 47564
rect 152595 47499 152661 47500
rect 152782 18869 152842 79731
rect 152963 76668 153029 76669
rect 152963 76604 152964 76668
rect 153028 76604 153029 76668
rect 152963 76603 153029 76604
rect 152779 18868 152845 18869
rect 152779 18804 152780 18868
rect 152844 18804 152845 18868
rect 152779 18803 152845 18804
rect 152966 13157 153026 76603
rect 153150 71229 153210 79731
rect 153883 78708 153949 78709
rect 153883 78644 153884 78708
rect 153948 78644 153949 78708
rect 153883 78643 153949 78644
rect 153147 71228 153213 71229
rect 153147 71164 153148 71228
rect 153212 71164 153213 71228
rect 153147 71163 153213 71164
rect 153886 40629 153946 78643
rect 154067 75852 154133 75853
rect 154067 75788 154068 75852
rect 154132 75788 154133 75852
rect 154067 75787 154133 75788
rect 153883 40628 153949 40629
rect 153883 40564 153884 40628
rect 153948 40564 153949 40628
rect 153883 40563 153949 40564
rect 154070 35189 154130 75787
rect 154067 35188 154133 35189
rect 154067 35124 154068 35188
rect 154132 35124 154133 35188
rect 154067 35123 154133 35124
rect 154254 16149 154314 79867
rect 154622 75989 154682 79867
rect 155358 78165 155418 79867
rect 155539 79660 155605 79661
rect 155539 79596 155540 79660
rect 155604 79596 155605 79660
rect 155539 79595 155605 79596
rect 155355 78164 155421 78165
rect 155355 78100 155356 78164
rect 155420 78100 155421 78164
rect 155355 78099 155421 78100
rect 154435 75988 154501 75989
rect 154435 75924 154436 75988
rect 154500 75924 154501 75988
rect 154435 75923 154501 75924
rect 154619 75988 154685 75989
rect 154619 75924 154620 75988
rect 154684 75924 154685 75988
rect 154619 75923 154685 75924
rect 154251 16148 154317 16149
rect 154251 16084 154252 16148
rect 154316 16084 154317 16148
rect 154251 16083 154317 16084
rect 154438 14789 154498 75923
rect 154794 48454 155414 78000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 14788 154501 14789
rect 154435 14724 154436 14788
rect 154500 14724 154501 14788
rect 154435 14723 154501 14724
rect 152963 13156 153029 13157
rect 152963 13092 152964 13156
rect 153028 13092 153029 13156
rect 152963 13091 153029 13092
rect 154794 12454 155414 47898
rect 155542 25533 155602 79595
rect 155723 76260 155789 76261
rect 155723 76196 155724 76260
rect 155788 76196 155789 76260
rect 155723 76195 155789 76196
rect 155539 25532 155605 25533
rect 155539 25468 155540 25532
rect 155604 25468 155605 25532
rect 155539 25467 155605 25468
rect 155726 16013 155786 76195
rect 156462 75989 156522 79867
rect 156643 79796 156709 79797
rect 156643 79732 156644 79796
rect 156708 79732 156709 79796
rect 156643 79731 156709 79732
rect 156459 75988 156525 75989
rect 156459 75924 156460 75988
rect 156524 75924 156525 75988
rect 156459 75923 156525 75924
rect 155723 16012 155789 16013
rect 155723 15948 155724 16012
rect 155788 15948 155789 16012
rect 155723 15947 155789 15948
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 151675 3636 151741 3637
rect 151675 3572 151676 3636
rect 151740 3572 151741 3636
rect 151675 3571 151741 3572
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 156646 8941 156706 79731
rect 156830 17373 156890 79867
rect 157011 77484 157077 77485
rect 157011 77420 157012 77484
rect 157076 77420 157077 77484
rect 157011 77419 157077 77420
rect 156827 17372 156893 17373
rect 156827 17308 156828 17372
rect 156892 17308 156893 17372
rect 156827 17307 156893 17308
rect 157014 14653 157074 77419
rect 157934 24173 157994 79867
rect 158483 79796 158549 79797
rect 158483 79732 158484 79796
rect 158548 79732 158549 79796
rect 158483 79731 158549 79732
rect 158299 78164 158365 78165
rect 158299 78100 158300 78164
rect 158364 78100 158365 78164
rect 158299 78099 158365 78100
rect 158115 78028 158181 78029
rect 158115 77964 158116 78028
rect 158180 77964 158181 78028
rect 158115 77963 158181 77964
rect 157931 24172 157997 24173
rect 157931 24108 157932 24172
rect 157996 24108 157997 24172
rect 157931 24107 157997 24108
rect 158118 18733 158178 77963
rect 158115 18732 158181 18733
rect 158115 18668 158116 18732
rect 158180 18668 158181 18732
rect 158115 18667 158181 18668
rect 158302 15877 158362 78099
rect 158299 15876 158365 15877
rect 158299 15812 158300 15876
rect 158364 15812 158365 15876
rect 158299 15811 158365 15812
rect 157011 14652 157077 14653
rect 157011 14588 157012 14652
rect 157076 14588 157077 14652
rect 157011 14587 157077 14588
rect 158486 11797 158546 79731
rect 158670 78573 158730 80139
rect 158851 79796 158917 79797
rect 158851 79732 158852 79796
rect 158916 79732 158917 79796
rect 158851 79731 158917 79732
rect 158667 78572 158733 78573
rect 158667 78508 158668 78572
rect 158732 78508 158733 78572
rect 158667 78507 158733 78508
rect 158854 21589 158914 79731
rect 159035 78708 159101 78709
rect 159035 78644 159036 78708
rect 159100 78644 159101 78708
rect 159035 78643 159101 78644
rect 158851 21588 158917 21589
rect 158851 21524 158852 21588
rect 158916 21524 158917 21588
rect 158851 21523 158917 21524
rect 158483 11796 158549 11797
rect 158483 11732 158484 11796
rect 158548 11732 158549 11796
rect 158483 11731 158549 11732
rect 156643 8940 156709 8941
rect 156643 8876 156644 8940
rect 156708 8876 156709 8940
rect 156643 8875 156709 8876
rect 159038 4997 159098 78643
rect 159774 78165 159834 80139
rect 160323 79932 160389 79933
rect 160323 79868 160324 79932
rect 160388 79868 160389 79932
rect 161059 79932 161125 79933
rect 161059 79930 161060 79932
rect 160323 79867 160389 79868
rect 160878 79870 161060 79930
rect 160326 78709 160386 79867
rect 160323 78708 160389 78709
rect 160323 78644 160324 78708
rect 160388 78644 160389 78708
rect 160323 78643 160389 78644
rect 160878 78570 160938 79870
rect 161059 79868 161060 79870
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 161795 79932 161861 79933
rect 161795 79868 161796 79932
rect 161860 79868 161861 79932
rect 161795 79867 161861 79868
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 162347 79932 162413 79933
rect 162347 79868 162348 79932
rect 162412 79868 162413 79932
rect 163451 79932 163517 79933
rect 163451 79930 163452 79932
rect 162347 79867 162413 79868
rect 163086 79870 163452 79930
rect 161798 78709 161858 79867
rect 161243 78708 161309 78709
rect 161243 78644 161244 78708
rect 161308 78644 161309 78708
rect 161243 78643 161309 78644
rect 161795 78708 161861 78709
rect 161795 78644 161796 78708
rect 161860 78644 161861 78708
rect 161795 78643 161861 78644
rect 160694 78510 160938 78570
rect 161059 78572 161125 78573
rect 159771 78164 159837 78165
rect 159771 78100 159772 78164
rect 159836 78100 159837 78164
rect 159771 78099 159837 78100
rect 159294 52954 159914 78000
rect 160694 61437 160754 78510
rect 161059 78508 161060 78572
rect 161124 78508 161125 78572
rect 161059 78507 161125 78508
rect 160875 78436 160941 78437
rect 160875 78372 160876 78436
rect 160940 78372 160941 78436
rect 160875 78371 160941 78372
rect 160691 61436 160757 61437
rect 160691 61372 160692 61436
rect 160756 61372 160757 61436
rect 160691 61371 160757 61372
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 160878 21453 160938 78371
rect 160875 21452 160941 21453
rect 160875 21388 160876 21452
rect 160940 21388 160941 21452
rect 160875 21387 160941 21388
rect 161062 20093 161122 78507
rect 161059 20092 161125 20093
rect 161059 20028 161060 20092
rect 161124 20028 161125 20092
rect 161059 20027 161125 20028
rect 161246 17237 161306 78643
rect 161982 77213 162042 79867
rect 162163 78708 162229 78709
rect 162163 78644 162164 78708
rect 162228 78644 162229 78708
rect 162163 78643 162229 78644
rect 161979 77212 162045 77213
rect 161979 77148 161980 77212
rect 162044 77148 162045 77212
rect 161979 77147 162045 77148
rect 162166 72725 162226 78643
rect 162163 72724 162229 72725
rect 162163 72660 162164 72724
rect 162228 72660 162229 72724
rect 162163 72659 162229 72660
rect 162350 21317 162410 79867
rect 162531 79660 162597 79661
rect 162531 79596 162532 79660
rect 162596 79596 162597 79660
rect 162531 79595 162597 79596
rect 162347 21316 162413 21317
rect 162347 21252 162348 21316
rect 162412 21252 162413 21316
rect 162347 21251 162413 21252
rect 161243 17236 161309 17237
rect 161243 17172 161244 17236
rect 161308 17172 161309 17236
rect 161243 17171 161309 17172
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 4996 159101 4997
rect 159035 4932 159036 4996
rect 159100 4932 159101 4996
rect 159035 4931 159101 4932
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 162534 14517 162594 79595
rect 162715 78708 162781 78709
rect 162715 78644 162716 78708
rect 162780 78644 162781 78708
rect 162715 78643 162781 78644
rect 162531 14516 162597 14517
rect 162531 14452 162532 14516
rect 162596 14452 162597 14516
rect 162531 14451 162597 14452
rect 162718 11661 162778 78643
rect 163086 77757 163146 79870
rect 163451 79868 163452 79870
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 164555 79932 164621 79933
rect 164555 79868 164556 79932
rect 164620 79868 164621 79932
rect 164555 79867 164621 79868
rect 163267 79660 163333 79661
rect 163267 79596 163268 79660
rect 163332 79596 163333 79660
rect 163267 79595 163333 79596
rect 163451 79660 163517 79661
rect 163451 79596 163452 79660
rect 163516 79596 163517 79660
rect 164187 79660 164253 79661
rect 164187 79658 164188 79660
rect 163451 79595 163517 79596
rect 163638 79598 164188 79658
rect 163083 77756 163149 77757
rect 163083 77692 163084 77756
rect 163148 77692 163149 77756
rect 163083 77691 163149 77692
rect 163270 77621 163330 79595
rect 163267 77620 163333 77621
rect 163267 77556 163268 77620
rect 163332 77556 163333 77620
rect 163267 77555 163333 77556
rect 163454 71093 163514 79595
rect 163451 71092 163517 71093
rect 163451 71028 163452 71092
rect 163516 71028 163517 71092
rect 163451 71027 163517 71028
rect 163638 19957 163698 79598
rect 164187 79596 164188 79598
rect 164252 79596 164253 79660
rect 164187 79595 164253 79596
rect 163794 57454 164414 78000
rect 164558 77621 164618 79867
rect 164923 78572 164989 78573
rect 164923 78508 164924 78572
rect 164988 78508 164989 78572
rect 164923 78507 164989 78508
rect 164555 77620 164621 77621
rect 164555 77556 164556 77620
rect 164620 77556 164621 77620
rect 164555 77555 164621 77556
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 19956 163701 19957
rect 163635 19892 163636 19956
rect 163700 19892 163701 19956
rect 163635 19891 163701 19892
rect 162715 11660 162781 11661
rect 162715 11596 162716 11660
rect 162780 11596 162781 11660
rect 162715 11595 162781 11596
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 10301 164986 78507
rect 165110 28253 165170 80139
rect 169523 80068 169589 80069
rect 169523 80004 169524 80068
rect 169588 80004 169589 80068
rect 169523 80003 169589 80004
rect 170811 80068 170877 80069
rect 170811 80004 170812 80068
rect 170876 80004 170877 80068
rect 170811 80003 170877 80004
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 166947 79932 167013 79933
rect 166947 79868 166948 79932
rect 167012 79930 167013 79932
rect 167315 79932 167381 79933
rect 167012 79870 167194 79930
rect 167012 79868 167013 79870
rect 166947 79867 167013 79868
rect 165107 28252 165173 28253
rect 165107 28188 165108 28252
rect 165172 28188 165173 28252
rect 165107 28187 165173 28188
rect 165294 27029 165354 79867
rect 165659 79796 165725 79797
rect 165659 79732 165660 79796
rect 165724 79732 165725 79796
rect 165659 79731 165725 79732
rect 165475 78844 165541 78845
rect 165475 78780 165476 78844
rect 165540 78780 165541 78844
rect 165475 78779 165541 78780
rect 165478 68237 165538 78779
rect 165662 78709 165722 79731
rect 165843 79660 165909 79661
rect 165843 79596 165844 79660
rect 165908 79596 165909 79660
rect 166763 79660 166829 79661
rect 166763 79658 166764 79660
rect 165843 79595 165909 79596
rect 166582 79598 166764 79658
rect 165846 78709 165906 79595
rect 165659 78708 165725 78709
rect 165659 78644 165660 78708
rect 165724 78644 165725 78708
rect 165659 78643 165725 78644
rect 165843 78708 165909 78709
rect 165843 78644 165844 78708
rect 165908 78644 165909 78708
rect 165843 78643 165909 78644
rect 166395 78708 166461 78709
rect 166395 78644 166396 78708
rect 166460 78644 166461 78708
rect 166395 78643 166461 78644
rect 165475 68236 165541 68237
rect 165475 68172 165476 68236
rect 165540 68172 165541 68236
rect 165475 68171 165541 68172
rect 166398 62933 166458 78643
rect 166395 62932 166461 62933
rect 166395 62868 166396 62932
rect 166460 62868 166461 62932
rect 166395 62867 166461 62868
rect 166582 32605 166642 79598
rect 166763 79596 166764 79598
rect 166828 79596 166829 79660
rect 166763 79595 166829 79596
rect 166763 77620 166829 77621
rect 166763 77556 166764 77620
rect 166828 77556 166829 77620
rect 166763 77555 166829 77556
rect 166579 32604 166645 32605
rect 166579 32540 166580 32604
rect 166644 32540 166645 32604
rect 166579 32539 166645 32540
rect 165291 27028 165357 27029
rect 165291 26964 165292 27028
rect 165356 26964 165357 27028
rect 165291 26963 165357 26964
rect 166766 13021 166826 77555
rect 167134 75173 167194 79870
rect 167315 79868 167316 79932
rect 167380 79868 167381 79932
rect 167315 79867 167381 79868
rect 167683 79932 167749 79933
rect 167683 79868 167684 79932
rect 167748 79868 167749 79932
rect 167683 79867 167749 79868
rect 167867 79932 167933 79933
rect 167867 79868 167868 79932
rect 167932 79868 167933 79932
rect 167867 79867 167933 79868
rect 168419 79932 168485 79933
rect 168419 79868 168420 79932
rect 168484 79868 168485 79932
rect 168419 79867 168485 79868
rect 168787 79932 168853 79933
rect 168787 79868 168788 79932
rect 168852 79868 168853 79932
rect 168787 79867 168853 79868
rect 169155 79932 169221 79933
rect 169155 79868 169156 79932
rect 169220 79868 169221 79932
rect 169155 79867 169221 79868
rect 167318 78165 167378 79867
rect 167686 78709 167746 79867
rect 167683 78708 167749 78709
rect 167683 78644 167684 78708
rect 167748 78644 167749 78708
rect 167683 78643 167749 78644
rect 167870 78573 167930 79867
rect 168051 79796 168117 79797
rect 168051 79732 168052 79796
rect 168116 79732 168117 79796
rect 168051 79731 168117 79732
rect 167867 78572 167933 78573
rect 167867 78508 167868 78572
rect 167932 78508 167933 78572
rect 167867 78507 167933 78508
rect 167315 78164 167381 78165
rect 167315 78100 167316 78164
rect 167380 78100 167381 78164
rect 167315 78099 167381 78100
rect 167683 78164 167749 78165
rect 167683 78100 167684 78164
rect 167748 78100 167749 78164
rect 167683 78099 167749 78100
rect 167131 75172 167197 75173
rect 167131 75108 167132 75172
rect 167196 75108 167197 75172
rect 167131 75107 167197 75108
rect 167686 30973 167746 78099
rect 168054 77890 168114 79731
rect 168422 78845 168482 79867
rect 168419 78844 168485 78845
rect 168419 78780 168420 78844
rect 168484 78780 168485 78844
rect 168419 78779 168485 78780
rect 168790 78165 168850 79867
rect 169158 78165 169218 79867
rect 169526 78573 169586 80003
rect 170075 79932 170141 79933
rect 170075 79868 170076 79932
rect 170140 79868 170141 79932
rect 170075 79867 170141 79868
rect 169891 79796 169957 79797
rect 169891 79732 169892 79796
rect 169956 79732 169957 79796
rect 169891 79731 169957 79732
rect 169523 78572 169589 78573
rect 169523 78508 169524 78572
rect 169588 78508 169589 78572
rect 169523 78507 169589 78508
rect 168787 78164 168853 78165
rect 168787 78100 168788 78164
rect 168852 78100 168853 78164
rect 168787 78099 168853 78100
rect 169155 78164 169221 78165
rect 169155 78100 169156 78164
rect 169220 78100 169221 78164
rect 169155 78099 169221 78100
rect 169523 78164 169589 78165
rect 169523 78100 169524 78164
rect 169588 78100 169589 78164
rect 169523 78099 169589 78100
rect 167870 77830 168114 77890
rect 167683 30972 167749 30973
rect 167683 30908 167684 30972
rect 167748 30908 167749 30972
rect 167683 30907 167749 30908
rect 167870 18597 167930 77830
rect 168051 77620 168117 77621
rect 168051 77556 168052 77620
rect 168116 77556 168117 77620
rect 168051 77555 168117 77556
rect 167867 18596 167933 18597
rect 167867 18532 167868 18596
rect 167932 18532 167933 18596
rect 167867 18531 167933 18532
rect 166763 13020 166829 13021
rect 166763 12956 166764 13020
rect 166828 12956 166829 13020
rect 166763 12955 166829 12956
rect 164923 10300 164989 10301
rect 164923 10236 164924 10300
rect 164988 10236 164989 10300
rect 164923 10235 164989 10236
rect 168054 4861 168114 77555
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169526 32469 169586 78099
rect 169894 76397 169954 79731
rect 170078 78709 170138 79867
rect 170443 79660 170509 79661
rect 170443 79596 170444 79660
rect 170508 79596 170509 79660
rect 170443 79595 170509 79596
rect 170446 78842 170506 79595
rect 170446 78782 170690 78842
rect 170075 78708 170141 78709
rect 170075 78644 170076 78708
rect 170140 78644 170141 78708
rect 170075 78643 170141 78644
rect 170443 78708 170509 78709
rect 170443 78644 170444 78708
rect 170508 78644 170509 78708
rect 170443 78643 170509 78644
rect 169891 76396 169957 76397
rect 169891 76332 169892 76396
rect 169956 76332 169957 76396
rect 169891 76331 169957 76332
rect 169523 32468 169589 32469
rect 169523 32404 169524 32468
rect 169588 32404 169589 32468
rect 169523 32403 169589 32404
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 4860 168117 4861
rect 168051 4796 168052 4860
rect 168116 4796 168117 4860
rect 168051 4795 168117 4796
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170446 21725 170506 78643
rect 170630 33829 170690 78782
rect 170627 33828 170693 33829
rect 170627 33764 170628 33828
rect 170692 33764 170693 33828
rect 170627 33763 170693 33764
rect 170814 26893 170874 80003
rect 171182 79933 171242 81091
rect 171915 81020 171981 81021
rect 171915 80956 171916 81020
rect 171980 80956 171981 81020
rect 171915 80955 171981 80956
rect 171363 80340 171429 80341
rect 171363 80276 171364 80340
rect 171428 80276 171429 80340
rect 171363 80275 171429 80276
rect 171547 80340 171613 80341
rect 171547 80276 171548 80340
rect 171612 80276 171613 80340
rect 171547 80275 171613 80276
rect 171179 79932 171245 79933
rect 171179 79868 171180 79932
rect 171244 79868 171245 79932
rect 171179 79867 171245 79868
rect 170995 79796 171061 79797
rect 170995 79732 170996 79796
rect 171060 79732 171061 79796
rect 170995 79731 171061 79732
rect 170998 78573 171058 79731
rect 170995 78572 171061 78573
rect 170995 78508 170996 78572
rect 171060 78508 171061 78572
rect 170995 78507 171061 78508
rect 171366 77893 171426 80275
rect 171550 78709 171610 80275
rect 171731 80204 171797 80205
rect 171731 80140 171732 80204
rect 171796 80140 171797 80204
rect 171731 80139 171797 80140
rect 171547 78708 171613 78709
rect 171547 78644 171548 78708
rect 171612 78644 171613 78708
rect 171547 78643 171613 78644
rect 171363 77892 171429 77893
rect 171363 77828 171364 77892
rect 171428 77828 171429 77892
rect 171363 77827 171429 77828
rect 170811 26892 170877 26893
rect 170811 26828 170812 26892
rect 170876 26828 170877 26892
rect 170811 26827 170877 26828
rect 170443 21724 170509 21725
rect 170443 21660 170444 21724
rect 170508 21660 170509 21724
rect 170443 21659 170509 21660
rect 171734 3501 171794 80139
rect 171918 79933 171978 80955
rect 172099 80748 172165 80749
rect 172099 80684 172100 80748
rect 172164 80684 172165 80748
rect 172099 80683 172165 80684
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 171915 79867 171981 79868
rect 172102 79797 172162 80683
rect 173019 80612 173085 80613
rect 173019 80548 173020 80612
rect 173084 80548 173085 80612
rect 173019 80547 173085 80548
rect 172835 80476 172901 80477
rect 172835 80412 172836 80476
rect 172900 80412 172901 80476
rect 172835 80411 172901 80412
rect 172838 80069 172898 80411
rect 173022 80069 173082 80547
rect 172835 80068 172901 80069
rect 172835 80004 172836 80068
rect 172900 80004 172901 80068
rect 172835 80003 172901 80004
rect 173019 80068 173085 80069
rect 173019 80004 173020 80068
rect 173084 80004 173085 80068
rect 173019 80003 173085 80004
rect 172283 79932 172349 79933
rect 172283 79868 172284 79932
rect 172348 79868 172349 79932
rect 172283 79867 172349 79868
rect 172467 79932 172533 79933
rect 172467 79868 172468 79932
rect 172532 79930 172533 79932
rect 172532 79870 173266 79930
rect 172532 79868 172533 79870
rect 172467 79867 172533 79868
rect 172099 79796 172165 79797
rect 172099 79732 172100 79796
rect 172164 79732 172165 79796
rect 172099 79731 172165 79732
rect 172099 78844 172165 78845
rect 172099 78780 172100 78844
rect 172164 78780 172165 78844
rect 172099 78779 172165 78780
rect 171915 75988 171981 75989
rect 171915 75924 171916 75988
rect 171980 75924 171981 75988
rect 171915 75923 171981 75924
rect 171731 3500 171797 3501
rect 171731 3436 171732 3500
rect 171796 3436 171797 3500
rect 171731 3435 171797 3436
rect 171918 3365 171978 75923
rect 172102 62797 172162 78779
rect 172286 77349 172346 79867
rect 172467 79796 172533 79797
rect 172467 79732 172468 79796
rect 172532 79732 172533 79796
rect 172467 79731 172533 79732
rect 172283 77348 172349 77349
rect 172283 77284 172284 77348
rect 172348 77284 172349 77348
rect 172283 77283 172349 77284
rect 172470 77213 172530 79731
rect 173206 78981 173266 79870
rect 173390 79117 173450 81227
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 173387 79116 173453 79117
rect 173387 79052 173388 79116
rect 173452 79052 173453 79116
rect 173387 79051 173453 79052
rect 173203 78980 173269 78981
rect 173203 78916 173204 78980
rect 173268 78916 173269 78980
rect 173203 78915 173269 78916
rect 172467 77212 172533 77213
rect 172467 77148 172468 77212
rect 172532 77148 172533 77212
rect 172467 77147 172533 77148
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172099 62796 172165 62797
rect 172099 62732 172100 62796
rect 172164 62732 172165 62796
rect 172099 62731 172165 62732
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 171915 3364 171981 3365
rect 171915 3300 171916 3364
rect 171980 3300 171981 3364
rect 171915 3299 171981 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 396582 78437 396642 696899
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 396579 78436 396645 78437
rect 396579 78372 396580 78436
rect 396644 78372 396645 78436
rect 396579 78371 396645 78372
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
