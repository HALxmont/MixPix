magic
tech sky130A
magscale 1 2
timestamp 1668297304
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 45278 700408 45284 700460
rect 45336 700448 45342 700460
rect 170306 700448 170312 700460
rect 45336 700420 170312 700448
rect 45336 700408 45342 700420
rect 170306 700408 170312 700420
rect 170364 700408 170370 700460
rect 364978 700408 364984 700460
rect 365036 700448 365042 700460
rect 397638 700448 397644 700460
rect 365036 700420 397644 700448
rect 365036 700408 365042 700420
rect 397638 700408 397644 700420
rect 397696 700408 397702 700460
rect 404998 700408 405004 700460
rect 405056 700448 405062 700460
rect 413646 700448 413652 700460
rect 405056 700420 413652 700448
rect 405056 700408 405062 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 44634 700340 44640 700392
rect 44692 700380 44698 700392
rect 235166 700380 235172 700392
rect 44692 700352 235172 700380
rect 44692 700340 44698 700352
rect 235166 700340 235172 700352
rect 235224 700340 235230 700392
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 293954 700380 293960 700392
rect 283892 700352 293960 700380
rect 283892 700340 283898 700352
rect 293954 700340 293960 700352
rect 294012 700340 294018 700392
rect 348786 700340 348792 700392
rect 348844 700380 348850 700392
rect 396442 700380 396448 700392
rect 348844 700352 396448 700380
rect 348844 700340 348850 700352
rect 396442 700340 396448 700352
rect 396500 700340 396506 700392
rect 403618 700340 403624 700392
rect 403676 700380 403682 700392
rect 478506 700380 478512 700392
rect 403676 700352 478512 700380
rect 403676 700340 403682 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 44726 700272 44732 700324
rect 44784 700312 44790 700324
rect 300118 700312 300124 700324
rect 44784 700284 300124 700312
rect 44784 700272 44790 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 397546 700312 397552 700324
rect 332560 700284 397552 700312
rect 332560 700272 332566 700284
rect 397546 700272 397552 700284
rect 397604 700272 397610 700324
rect 400858 700272 400864 700324
rect 400916 700312 400922 700324
rect 543458 700312 543464 700324
rect 400916 700284 543464 700312
rect 400916 700272 400922 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 198734 699660 198740 699712
rect 198792 699700 198798 699712
rect 202782 699700 202788 699712
rect 198792 699672 202788 699700
rect 198792 699660 198798 699672
rect 202782 699660 202788 699672
rect 202840 699660 202846 699712
rect 258718 699660 258724 699712
rect 258776 699700 258782 699712
rect 267642 699700 267648 699712
rect 258776 699672 267648 699700
rect 258776 699660 258782 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 398098 696940 398104 696992
rect 398156 696980 398162 696992
rect 580166 696980 580172 696992
rect 398156 696952 580172 696980
rect 398156 696940 398162 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 187970 694764 187976 694816
rect 188028 694804 188034 694816
rect 198734 694804 198740 694816
rect 188028 694776 198740 694804
rect 188028 694764 188034 694776
rect 198734 694764 198740 694776
rect 198792 694764 198798 694816
rect 293954 693404 293960 693456
rect 294012 693444 294018 693456
rect 305638 693444 305644 693456
rect 294012 693416 305644 693444
rect 294012 693404 294018 693416
rect 305638 693404 305644 693416
rect 305696 693404 305702 693456
rect 185578 691364 185584 691416
rect 185636 691404 185642 691416
rect 187970 691404 187976 691416
rect 185636 691376 187976 691404
rect 185636 691364 185642 691376
rect 187970 691364 187976 691376
rect 188028 691364 188034 691416
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 399478 683136 399484 683188
rect 399536 683176 399542 683188
rect 580166 683176 580172 683188
rect 399536 683148 580172 683176
rect 399536 683136 399542 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 253934 681776 253940 681828
rect 253992 681816 253998 681828
rect 258718 681816 258724 681828
rect 253992 681788 258724 681816
rect 253992 681776 253998 681788
rect 258718 681776 258724 681788
rect 258776 681776 258782 681828
rect 305638 679600 305644 679652
rect 305696 679640 305702 679652
rect 322198 679640 322204 679652
rect 305696 679612 322204 679640
rect 305696 679600 305702 679612
rect 322198 679600 322204 679612
rect 322256 679600 322262 679652
rect 239398 678240 239404 678292
rect 239456 678280 239462 678292
rect 253934 678280 253940 678292
rect 239456 678252 253940 678280
rect 239456 678240 239462 678252
rect 253934 678240 253940 678252
rect 253992 678240 253998 678292
rect 147766 678036 147772 678088
rect 147824 678076 147830 678088
rect 153194 678076 153200 678088
rect 147824 678048 153200 678076
rect 147824 678036 147830 678048
rect 153194 678036 153200 678048
rect 153252 678036 153258 678088
rect 147030 675520 147036 675572
rect 147088 675560 147094 675572
rect 147766 675560 147772 675572
rect 147088 675532 147772 675560
rect 147088 675520 147094 675532
rect 147766 675520 147772 675532
rect 147824 675520 147830 675572
rect 236638 671168 236644 671220
rect 236696 671208 236702 671220
rect 239398 671208 239404 671220
rect 236696 671180 239404 671208
rect 236696 671168 236702 671180
rect 239398 671168 239404 671180
rect 239456 671168 239462 671220
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 18598 670732 18604 670744
rect 3568 670704 18604 670732
rect 3568 670692 3574 670704
rect 18598 670692 18604 670704
rect 18656 670692 18662 670744
rect 145558 667836 145564 667888
rect 145616 667876 145622 667888
rect 147030 667876 147036 667888
rect 145616 667848 147036 667876
rect 145616 667836 145622 667848
rect 147030 667836 147036 667848
rect 147088 667836 147094 667888
rect 231302 662396 231308 662448
rect 231360 662436 231366 662448
rect 236638 662436 236644 662448
rect 231360 662408 236644 662436
rect 231360 662396 231366 662408
rect 236638 662396 236644 662408
rect 236696 662396 236702 662448
rect 224218 659744 224224 659796
rect 224276 659784 224282 659796
rect 231302 659784 231308 659796
rect 224276 659756 231308 659784
rect 224276 659744 224282 659756
rect 231302 659744 231308 659756
rect 231360 659744 231366 659796
rect 142798 657976 142804 658028
rect 142856 658016 142862 658028
rect 145558 658016 145564 658028
rect 142856 657988 145564 658016
rect 142856 657976 142862 657988
rect 145558 657976 145564 657988
rect 145616 657976 145622 658028
rect 177850 653352 177856 653404
rect 177908 653392 177914 653404
rect 185578 653392 185584 653404
rect 177908 653364 185584 653392
rect 177908 653352 177914 653364
rect 185578 653352 185584 653364
rect 185636 653352 185642 653404
rect 142798 652780 142804 652792
rect 139412 652752 142804 652780
rect 138382 652672 138388 652724
rect 138440 652712 138446 652724
rect 139412 652712 139440 652752
rect 142798 652740 142804 652752
rect 142856 652740 142862 652792
rect 138440 652684 139440 652712
rect 138440 652672 138446 652684
rect 174814 646688 174820 646740
rect 174872 646728 174878 646740
rect 177850 646728 177856 646740
rect 174872 646700 177856 646728
rect 174872 646688 174878 646700
rect 177850 646688 177856 646700
rect 177908 646688 177914 646740
rect 138382 644484 138388 644496
rect 136652 644456 138388 644484
rect 135898 644376 135904 644428
rect 135956 644416 135962 644428
rect 136652 644416 136680 644456
rect 138382 644444 138388 644456
rect 138440 644444 138446 644496
rect 135956 644388 136680 644416
rect 135956 644376 135962 644388
rect 396718 643084 396724 643136
rect 396776 643124 396782 643136
rect 580166 643124 580172 643136
rect 396776 643096 580172 643124
rect 396776 643084 396782 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 214558 638868 214564 638920
rect 214616 638908 214622 638920
rect 218054 638908 218060 638920
rect 214616 638880 218060 638908
rect 214616 638868 214622 638880
rect 218054 638868 218060 638880
rect 218112 638868 218118 638920
rect 152458 638188 152464 638240
rect 152516 638228 152522 638240
rect 174814 638228 174820 638240
rect 152516 638200 174820 638228
rect 152516 638188 152522 638200
rect 174814 638188 174820 638200
rect 174872 638188 174878 638240
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 7558 632108 7564 632120
rect 3568 632080 7564 632108
rect 3568 632068 3574 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 210418 632068 210424 632120
rect 210476 632108 210482 632120
rect 214558 632108 214564 632120
rect 210476 632080 214564 632108
rect 210476 632068 210482 632080
rect 214558 632068 214564 632080
rect 214616 632068 214622 632120
rect 133138 630640 133144 630692
rect 133196 630680 133202 630692
rect 135898 630680 135904 630692
rect 133196 630652 135904 630680
rect 133196 630640 133202 630652
rect 135898 630640 135904 630652
rect 135956 630640 135962 630692
rect 417418 630640 417424 630692
rect 417476 630680 417482 630692
rect 579982 630680 579988 630692
rect 417476 630652 579988 630680
rect 417476 630640 417482 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 129734 623772 129740 623824
rect 129792 623812 129798 623824
rect 133138 623812 133144 623824
rect 129792 623784 133144 623812
rect 129792 623772 129798 623784
rect 133138 623772 133144 623784
rect 133196 623772 133202 623824
rect 214558 623024 214564 623076
rect 214616 623064 214622 623076
rect 224218 623064 224224 623076
rect 214616 623036 224224 623064
rect 214616 623024 214622 623036
rect 224218 623024 224224 623036
rect 224276 623024 224282 623076
rect 322198 622412 322204 622464
rect 322256 622452 322262 622464
rect 324958 622452 324964 622464
rect 322256 622424 324964 622452
rect 322256 622412 322262 622424
rect 324958 622412 324964 622424
rect 325016 622412 325022 622464
rect 128998 620984 129004 621036
rect 129056 621024 129062 621036
rect 129734 621024 129740 621036
rect 129056 620996 129740 621024
rect 129056 620984 129062 620996
rect 129734 620984 129740 620996
rect 129792 620984 129798 621036
rect 196618 620236 196624 620288
rect 196676 620276 196682 620288
rect 214558 620276 214564 620288
rect 196676 620248 214564 620276
rect 196676 620236 196682 620248
rect 214558 620236 214564 620248
rect 214616 620236 214622 620288
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 21358 618304 21364 618316
rect 3568 618276 21364 618304
rect 3568 618264 3574 618276
rect 21358 618264 21364 618276
rect 21416 618264 21422 618316
rect 207014 611872 207020 611924
rect 207072 611912 207078 611924
rect 210418 611912 210424 611924
rect 207072 611884 210424 611912
rect 207072 611872 207078 611884
rect 210418 611872 210424 611884
rect 210476 611872 210482 611924
rect 130378 609220 130384 609272
rect 130436 609260 130442 609272
rect 207014 609260 207020 609272
rect 130436 609232 207020 609260
rect 130436 609220 130442 609232
rect 207014 609220 207020 609232
rect 207072 609220 207078 609272
rect 189074 605072 189080 605124
rect 189132 605112 189138 605124
rect 196618 605112 196624 605124
rect 189132 605084 196624 605112
rect 189132 605072 189138 605084
rect 196618 605072 196624 605084
rect 196676 605072 196682 605124
rect 181438 600448 181444 600500
rect 181496 600488 181502 600500
rect 189074 600488 189080 600500
rect 181496 600460 189080 600488
rect 181496 600448 181502 600460
rect 189074 600448 189080 600460
rect 189132 600448 189138 600500
rect 127618 598816 127624 598868
rect 127676 598856 127682 598868
rect 130378 598856 130384 598868
rect 127676 598828 130384 598856
rect 127676 598816 127682 598828
rect 130378 598816 130384 598828
rect 130436 598816 130442 598868
rect 149330 594804 149336 594856
rect 149388 594844 149394 594856
rect 152458 594844 152464 594856
rect 149388 594816 152464 594844
rect 149388 594804 149394 594816
rect 152458 594804 152464 594816
rect 152516 594804 152522 594856
rect 146938 592016 146944 592068
rect 146996 592056 147002 592068
rect 149330 592056 149336 592068
rect 146996 592028 149336 592056
rect 146996 592016 147002 592028
rect 149330 592016 149336 592028
rect 149388 592016 149394 592068
rect 159358 589908 159364 589960
rect 159416 589948 159422 589960
rect 181438 589948 181444 589960
rect 159416 589920 181444 589948
rect 159416 589908 159422 589920
rect 181438 589908 181444 589920
rect 181496 589908 181502 589960
rect 124858 581612 124864 581664
rect 124916 581652 124922 581664
rect 127618 581652 127624 581664
rect 124916 581624 127624 581652
rect 124916 581612 124922 581624
rect 127618 581612 127624 581624
rect 127676 581612 127682 581664
rect 2774 579912 2780 579964
rect 2832 579952 2838 579964
rect 4890 579952 4896 579964
rect 2832 579924 4896 579952
rect 2832 579912 2838 579924
rect 4890 579912 4896 579924
rect 4948 579912 4954 579964
rect 414658 576852 414664 576904
rect 414716 576892 414722 576904
rect 580166 576892 580172 576904
rect 414716 576864 580172 576892
rect 414716 576852 414722 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 324958 570596 324964 570648
rect 325016 570636 325022 570648
rect 329098 570636 329104 570648
rect 325016 570608 329104 570636
rect 325016 570596 325022 570608
rect 329098 570596 329104 570608
rect 329156 570596 329162 570648
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 31018 565876 31024 565888
rect 3108 565848 31024 565876
rect 3108 565836 3114 565848
rect 31018 565836 31024 565848
rect 31076 565836 31082 565888
rect 141418 565088 141424 565140
rect 141476 565128 141482 565140
rect 146938 565128 146944 565140
rect 141476 565100 146944 565128
rect 141476 565088 141482 565100
rect 146938 565088 146944 565100
rect 146996 565088 147002 565140
rect 138014 554752 138020 554804
rect 138072 554792 138078 554804
rect 141418 554792 141424 554804
rect 138072 554764 141424 554792
rect 138072 554752 138078 554764
rect 141418 554752 141424 554764
rect 141476 554752 141482 554804
rect 135898 550536 135904 550588
rect 135956 550576 135962 550588
rect 138014 550576 138020 550588
rect 135956 550548 138020 550576
rect 135956 550536 135962 550548
rect 138014 550536 138020 550548
rect 138072 550536 138078 550588
rect 155218 542512 155224 542564
rect 155276 542552 155282 542564
rect 159358 542552 159364 542564
rect 155276 542524 159364 542552
rect 155276 542512 155282 542524
rect 159358 542512 159364 542524
rect 159416 542512 159422 542564
rect 127618 540880 127624 540932
rect 127676 540920 127682 540932
rect 128998 540920 129004 540932
rect 127676 540892 129004 540920
rect 127676 540880 127682 540892
rect 128998 540880 129004 540892
rect 129056 540880 129062 540932
rect 329098 532652 329104 532704
rect 329156 532692 329162 532704
rect 331214 532692 331220 532704
rect 329156 532664 331220 532692
rect 329156 532652 329162 532664
rect 331214 532652 331220 532664
rect 331272 532652 331278 532704
rect 126238 529864 126244 529916
rect 126296 529904 126302 529916
rect 127618 529904 127624 529916
rect 126296 529876 127624 529904
rect 126296 529864 126302 529876
rect 127618 529864 127624 529876
rect 127676 529864 127682 529916
rect 331214 529184 331220 529236
rect 331272 529224 331278 529236
rect 341518 529224 341524 529236
rect 331272 529196 341524 529224
rect 331272 529184 331278 529196
rect 341518 529184 341524 529196
rect 341576 529184 341582 529236
rect 3510 527824 3516 527876
rect 3568 527864 3574 527876
rect 8938 527864 8944 527876
rect 3568 527836 8944 527864
rect 3568 527824 3574 527836
rect 8938 527824 8944 527836
rect 8996 527824 9002 527876
rect 413278 524424 413284 524476
rect 413336 524464 413342 524476
rect 580074 524464 580080 524476
rect 413336 524436 580080 524464
rect 413336 524424 413342 524436
rect 580074 524424 580080 524436
rect 580132 524424 580138 524476
rect 124214 520208 124220 520260
rect 124272 520248 124278 520260
rect 126238 520248 126244 520260
rect 124272 520220 126244 520248
rect 124272 520208 124278 520220
rect 126238 520208 126244 520220
rect 126296 520208 126302 520260
rect 122098 518916 122104 518968
rect 122156 518956 122162 518968
rect 124858 518956 124864 518968
rect 122156 518928 124864 518956
rect 122156 518916 122162 518928
rect 124858 518916 124864 518928
rect 124916 518916 124922 518968
rect 341518 517896 341524 517948
rect 341576 517936 341582 517948
rect 343634 517936 343640 517948
rect 341576 517908 343640 517936
rect 341576 517896 341582 517908
rect 343634 517896 343640 517908
rect 343692 517896 343698 517948
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 32398 514808 32404 514820
rect 3568 514780 32404 514808
rect 3568 514768 3574 514780
rect 32398 514768 32404 514780
rect 32456 514768 32462 514820
rect 123478 514768 123484 514820
rect 123536 514808 123542 514820
rect 124214 514808 124220 514820
rect 123536 514780 124220 514808
rect 123536 514768 123542 514780
rect 124214 514768 124220 514780
rect 124272 514768 124278 514820
rect 343634 513272 343640 513324
rect 343692 513312 343698 513324
rect 347038 513312 347044 513324
rect 343692 513284 347044 513312
rect 343692 513272 343698 513284
rect 347038 513272 347044 513284
rect 347096 513272 347102 513324
rect 118970 511844 118976 511896
rect 119028 511884 119034 511896
rect 122098 511884 122104 511896
rect 119028 511856 122104 511884
rect 119028 511844 119034 511856
rect 122098 511844 122104 511856
rect 122156 511844 122162 511896
rect 116026 507832 116032 507884
rect 116084 507872 116090 507884
rect 118970 507872 118976 507884
rect 116084 507844 118976 507872
rect 116084 507832 116090 507844
rect 118970 507832 118976 507844
rect 119028 507832 119034 507884
rect 102778 502936 102784 502988
rect 102836 502976 102842 502988
rect 116026 502976 116032 502988
rect 102836 502948 116032 502976
rect 102836 502936 102842 502948
rect 116026 502936 116032 502948
rect 116084 502936 116090 502988
rect 100018 498176 100024 498228
rect 100076 498216 100082 498228
rect 102778 498216 102784 498228
rect 100076 498188 102784 498216
rect 100076 498176 100082 498188
rect 102778 498176 102784 498188
rect 102836 498176 102842 498228
rect 152458 480292 152464 480344
rect 152516 480332 152522 480344
rect 155218 480332 155224 480344
rect 152516 480304 155224 480332
rect 152516 480292 152522 480304
rect 155218 480292 155224 480304
rect 155276 480292 155282 480344
rect 347038 476008 347044 476060
rect 347096 476048 347102 476060
rect 353294 476048 353300 476060
rect 347096 476020 353300 476048
rect 347096 476008 347102 476020
rect 353294 476008 353300 476020
rect 353352 476008 353358 476060
rect 3510 474716 3516 474768
rect 3568 474756 3574 474768
rect 13078 474756 13084 474768
rect 3568 474728 13084 474756
rect 3568 474716 3574 474728
rect 13078 474716 13084 474728
rect 13136 474716 13142 474768
rect 353294 472404 353300 472456
rect 353352 472444 353358 472456
rect 356054 472444 356060 472456
rect 353352 472416 356060 472444
rect 353352 472404 353358 472416
rect 356054 472404 356060 472416
rect 356112 472404 356118 472456
rect 522298 470568 522304 470620
rect 522356 470608 522362 470620
rect 580074 470608 580080 470620
rect 522356 470580 580080 470608
rect 522356 470568 522362 470580
rect 580074 470568 580080 470580
rect 580132 470568 580138 470620
rect 142798 468460 142804 468512
rect 142856 468500 142862 468512
rect 152458 468500 152464 468512
rect 142856 468472 152464 468500
rect 142856 468460 142862 468472
rect 152458 468460 152464 468472
rect 152516 468460 152522 468512
rect 356054 467712 356060 467764
rect 356112 467752 356118 467764
rect 358998 467752 359004 467764
rect 356112 467724 359004 467752
rect 356112 467712 356118 467724
rect 358998 467712 359004 467724
rect 359056 467712 359062 467764
rect 97258 464720 97264 464772
rect 97316 464760 97322 464772
rect 100018 464760 100024 464772
rect 97316 464732 100024 464760
rect 97316 464720 97322 464732
rect 100018 464720 100024 464732
rect 100076 464720 100082 464772
rect 358998 464312 359004 464364
rect 359056 464352 359062 464364
rect 370498 464352 370504 464364
rect 359056 464324 370504 464352
rect 359056 464312 359062 464324
rect 370498 464312 370504 464324
rect 370556 464312 370562 464364
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 22738 462380 22744 462392
rect 3568 462352 22744 462380
rect 3568 462340 3574 462352
rect 22738 462340 22744 462352
rect 22796 462340 22802 462392
rect 370498 459484 370504 459536
rect 370556 459524 370562 459536
rect 376294 459524 376300 459536
rect 370556 459496 376300 459524
rect 370556 459484 370562 459496
rect 376294 459484 376300 459496
rect 376352 459484 376358 459536
rect 88978 458804 88984 458856
rect 89036 458844 89042 458856
rect 97258 458844 97264 458856
rect 89036 458816 97264 458844
rect 89036 458804 89042 458816
rect 97258 458804 97264 458816
rect 97316 458804 97322 458856
rect 376294 456356 376300 456408
rect 376352 456396 376358 456408
rect 381538 456396 381544 456408
rect 376352 456368 381544 456396
rect 376352 456356 376358 456368
rect 381538 456356 381544 456368
rect 381596 456356 381602 456408
rect 120718 453296 120724 453348
rect 120776 453336 120782 453348
rect 142798 453336 142804 453348
rect 120776 453308 142804 453336
rect 120776 453296 120782 453308
rect 142798 453296 142804 453308
rect 142856 453296 142862 453348
rect 381538 437384 381544 437436
rect 381596 437424 381602 437436
rect 384298 437424 384304 437436
rect 381596 437396 384304 437424
rect 381596 437384 381602 437396
rect 384298 437384 384304 437396
rect 384356 437384 384362 437436
rect 125502 425688 125508 425740
rect 125560 425728 125566 425740
rect 135898 425728 135904 425740
rect 125560 425700 135904 425728
rect 125560 425688 125566 425700
rect 135898 425688 135904 425700
rect 135956 425688 135962 425740
rect 113818 422900 113824 422952
rect 113876 422940 113882 422952
rect 125502 422940 125508 422952
rect 113876 422912 125508 422940
rect 113876 422900 113882 422912
rect 125502 422900 125508 422912
rect 125560 422900 125566 422952
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 10318 422328 10324 422340
rect 3384 422300 10324 422328
rect 3384 422288 3390 422300
rect 10318 422288 10324 422300
rect 10376 422288 10382 422340
rect 122098 420180 122104 420232
rect 122156 420220 122162 420232
rect 123478 420220 123484 420232
rect 122156 420192 123484 420220
rect 122156 420180 122162 420192
rect 123478 420180 123484 420192
rect 123536 420180 123542 420232
rect 86218 419500 86224 419552
rect 86276 419540 86282 419552
rect 88978 419540 88984 419552
rect 86276 419512 88984 419540
rect 86276 419500 86282 419512
rect 88978 419500 88984 419512
rect 89036 419500 89042 419552
rect 409138 418140 409144 418192
rect 409196 418180 409202 418192
rect 580074 418180 580080 418192
rect 409196 418152 580080 418180
rect 409196 418140 409202 418152
rect 580074 418140 580080 418152
rect 580132 418140 580138 418192
rect 384298 415352 384304 415404
rect 384356 415392 384362 415404
rect 387702 415392 387708 415404
rect 384356 415364 387708 415392
rect 384356 415352 384362 415364
rect 387702 415352 387708 415364
rect 387760 415352 387766 415404
rect 387702 411884 387708 411936
rect 387760 411924 387766 411936
rect 396534 411924 396540 411936
rect 387760 411896 396540 411924
rect 387760 411884 387766 411896
rect 396534 411884 396540 411896
rect 396592 411884 396598 411936
rect 83458 410116 83464 410168
rect 83516 410156 83522 410168
rect 86218 410156 86224 410168
rect 83516 410128 86224 410156
rect 83516 410116 83522 410128
rect 86218 410116 86224 410128
rect 86276 410116 86282 410168
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 28258 409884 28264 409896
rect 3384 409856 28264 409884
rect 3384 409844 3390 409856
rect 28258 409844 28264 409856
rect 28316 409844 28322 409896
rect 396810 404336 396816 404388
rect 396868 404376 396874 404388
rect 580074 404376 580080 404388
rect 396868 404348 580080 404376
rect 396868 404336 396874 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 119338 401616 119344 401668
rect 119396 401656 119402 401668
rect 122098 401656 122104 401668
rect 119396 401628 122104 401656
rect 119396 401616 119402 401628
rect 122098 401616 122104 401628
rect 122156 401616 122162 401668
rect 116578 398828 116584 398880
rect 116636 398868 116642 398880
rect 119338 398868 119344 398880
rect 116636 398840 119344 398868
rect 116636 398828 116642 398840
rect 119338 398828 119344 398840
rect 119396 398828 119402 398880
rect 69658 396720 69664 396772
rect 69716 396760 69722 396772
rect 136634 396760 136640 396772
rect 69716 396732 136640 396760
rect 69716 396720 69722 396732
rect 136634 396720 136640 396732
rect 136692 396720 136698 396772
rect 68278 384956 68284 385008
rect 68336 384996 68342 385008
rect 69658 384996 69664 385008
rect 68336 384968 69664 384996
rect 68336 384956 68342 384968
rect 69658 384956 69664 384968
rect 69716 384956 69722 385008
rect 102042 384276 102048 384328
rect 102100 384316 102106 384328
rect 113818 384316 113824 384328
rect 102100 384288 113824 384316
rect 102100 384276 102106 384288
rect 113818 384276 113824 384288
rect 113876 384276 113882 384328
rect 398190 378156 398196 378208
rect 398248 378196 398254 378208
rect 580074 378196 580080 378208
rect 398248 378168 580080 378196
rect 398248 378156 398254 378168
rect 580074 378156 580080 378168
rect 580132 378156 580138 378208
rect 98638 377748 98644 377800
rect 98696 377788 98702 377800
rect 102042 377788 102048 377800
rect 98696 377760 102048 377788
rect 98696 377748 98702 377760
rect 102042 377748 102048 377760
rect 102100 377748 102106 377800
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 14458 371260 14464 371272
rect 3384 371232 14464 371260
rect 3384 371220 3390 371232
rect 14458 371220 14464 371232
rect 14516 371220 14522 371272
rect 77938 371220 77944 371272
rect 77996 371260 78002 371272
rect 83458 371260 83464 371272
rect 77996 371232 83464 371260
rect 77996 371220 78002 371232
rect 83458 371220 83464 371232
rect 83516 371220 83522 371272
rect 114922 370744 114928 370796
rect 114980 370784 114986 370796
rect 116578 370784 116584 370796
rect 114980 370756 116584 370784
rect 114980 370744 114986 370756
rect 116578 370744 116584 370756
rect 116636 370744 116642 370796
rect 112438 367752 112444 367804
rect 112496 367792 112502 367804
rect 114922 367792 114928 367804
rect 112496 367764 114928 367792
rect 112496 367752 112502 367764
rect 114922 367752 114928 367764
rect 114980 367752 114986 367804
rect 418798 364352 418804 364404
rect 418856 364392 418862 364404
rect 579798 364392 579804 364404
rect 418856 364364 579804 364392
rect 418856 364352 418862 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 117314 362924 117320 362976
rect 117372 362964 117378 362976
rect 120718 362964 120724 362976
rect 117372 362936 120724 362964
rect 117372 362924 117378 362936
rect 120718 362924 120724 362936
rect 120776 362924 120782 362976
rect 65426 358776 65432 358828
rect 65484 358816 65490 358828
rect 68278 358816 68284 358828
rect 65484 358788 68284 358816
rect 65484 358776 65490 358788
rect 68278 358776 68284 358788
rect 68336 358776 68342 358828
rect 64138 358096 64144 358148
rect 64196 358136 64202 358148
rect 65426 358136 65432 358148
rect 64196 358108 65432 358136
rect 64196 358096 64202 358108
rect 65426 358096 65432 358108
rect 65484 358096 65490 358148
rect 92474 358028 92480 358080
rect 92532 358068 92538 358080
rect 98638 358068 98644 358080
rect 92532 358040 98644 358068
rect 92532 358028 92538 358040
rect 98638 358028 98644 358040
rect 98696 358028 98702 358080
rect 113174 357008 113180 357060
rect 113232 357048 113238 357060
rect 117314 357048 117320 357060
rect 113232 357020 117320 357048
rect 113232 357008 113238 357020
rect 117314 357008 117320 357020
rect 117372 357008 117378 357060
rect 79318 355308 79324 355360
rect 79376 355348 79382 355360
rect 92474 355348 92480 355360
rect 79376 355320 92480 355348
rect 79376 355308 79382 355320
rect 92474 355308 92480 355320
rect 92532 355308 92538 355360
rect 111058 353268 111064 353320
rect 111116 353308 111122 353320
rect 112438 353308 112444 353320
rect 111116 353280 112444 353308
rect 111116 353268 111122 353280
rect 112438 353268 112444 353280
rect 112496 353268 112502 353320
rect 396902 351908 396908 351960
rect 396960 351948 396966 351960
rect 580074 351948 580080 351960
rect 396960 351920 580080 351948
rect 396960 351908 396966 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 45830 349800 45836 349852
rect 45888 349840 45894 349852
rect 77938 349840 77944 349852
rect 45888 349812 77944 349840
rect 45888 349800 45894 349812
rect 77938 349800 77944 349812
rect 77996 349800 78002 349852
rect 106918 348712 106924 348764
rect 106976 348752 106982 348764
rect 113174 348752 113180 348764
rect 106976 348724 113180 348752
rect 106976 348712 106982 348724
rect 113174 348712 113180 348724
rect 113232 348712 113238 348764
rect 109770 343612 109776 343664
rect 109828 343652 109834 343664
rect 111058 343652 111064 343664
rect 109828 343624 111064 343652
rect 109828 343612 109834 343624
rect 111058 343612 111064 343624
rect 111116 343612 111122 343664
rect 108298 340008 108304 340060
rect 108356 340048 108362 340060
rect 109770 340048 109776 340060
rect 108356 340020 109776 340048
rect 108356 340008 108362 340020
rect 109770 340008 109776 340020
rect 109828 340008 109834 340060
rect 104526 338240 104532 338292
rect 104584 338280 104590 338292
rect 106918 338280 106924 338292
rect 104584 338252 106924 338280
rect 104584 338240 104590 338252
rect 106918 338240 106924 338252
rect 106976 338240 106982 338292
rect 100754 335316 100760 335368
rect 100812 335356 100818 335368
rect 104526 335356 104532 335368
rect 100812 335328 104532 335356
rect 100812 335316 100818 335328
rect 104526 335316 104532 335328
rect 104584 335316 104590 335368
rect 76558 333208 76564 333260
rect 76616 333248 76622 333260
rect 100754 333248 100760 333260
rect 76616 333220 100760 333248
rect 76616 333208 76622 333220
rect 100754 333208 100760 333220
rect 100812 333208 100818 333260
rect 76650 329536 76656 329588
rect 76708 329576 76714 329588
rect 79318 329576 79324 329588
rect 76708 329548 79324 329576
rect 76708 329536 76714 329548
rect 79318 329536 79324 329548
rect 79376 329536 79382 329588
rect 72418 321376 72424 321428
rect 72476 321416 72482 321428
rect 76558 321416 76564 321428
rect 72476 321388 76564 321416
rect 72476 321376 72482 321388
rect 76558 321376 76564 321388
rect 76616 321376 76622 321428
rect 62758 319404 62764 319456
rect 62816 319444 62822 319456
rect 64138 319444 64144 319456
rect 62816 319416 64144 319444
rect 62816 319404 62822 319416
rect 64138 319404 64144 319416
rect 64196 319404 64202 319456
rect 73798 318996 73804 319048
rect 73856 319036 73862 319048
rect 76650 319036 76656 319048
rect 73856 319008 76656 319036
rect 73856 318996 73862 319008
rect 76650 318996 76656 319008
rect 76708 318996 76714 319048
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 26878 318832 26884 318844
rect 3200 318804 26884 318832
rect 3200 318792 3206 318804
rect 26878 318792 26884 318804
rect 26936 318792 26942 318844
rect 58618 315256 58624 315308
rect 58676 315296 58682 315308
rect 72418 315296 72424 315308
rect 58676 315268 72424 315296
rect 58676 315256 58682 315268
rect 72418 315256 72424 315268
rect 72476 315256 72482 315308
rect 407758 311856 407764 311908
rect 407816 311896 407822 311908
rect 579982 311896 579988 311908
rect 407816 311868 579988 311896
rect 407816 311856 407822 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 62850 305600 62856 305652
rect 62908 305640 62914 305652
rect 108298 305640 108304 305652
rect 62908 305612 108304 305640
rect 62908 305600 62914 305612
rect 108298 305600 108304 305612
rect 108356 305600 108362 305652
rect 61470 299412 61476 299464
rect 61528 299452 61534 299464
rect 62758 299452 62764 299464
rect 61528 299424 62764 299452
rect 61528 299412 61534 299424
rect 62758 299412 62764 299424
rect 62816 299412 62822 299464
rect 54478 298732 54484 298784
rect 54536 298772 54542 298784
rect 58618 298772 58624 298784
rect 54536 298744 58624 298772
rect 54536 298732 54542 298744
rect 58618 298732 58624 298744
rect 58676 298732 58682 298784
rect 396994 298120 397000 298172
rect 397052 298160 397058 298172
rect 579982 298160 579988 298172
rect 397052 298132 579988 298160
rect 397052 298120 397058 298132
rect 579982 298120 579988 298132
rect 580040 298120 580046 298172
rect 68278 295332 68284 295384
rect 68336 295372 68342 295384
rect 73798 295372 73804 295384
rect 68336 295344 73804 295372
rect 68336 295332 68342 295344
rect 73798 295332 73804 295344
rect 73856 295332 73862 295384
rect 61194 294040 61200 294092
rect 61252 294080 61258 294092
rect 62850 294080 62856 294092
rect 61252 294052 62856 294080
rect 61252 294040 61258 294052
rect 62850 294040 62856 294052
rect 62908 294040 62914 294092
rect 59998 293972 60004 294024
rect 60056 294012 60062 294024
rect 61470 294012 61476 294024
rect 60056 293984 61476 294012
rect 60056 293972 60062 293984
rect 61470 293972 61476 293984
rect 61528 293972 61534 294024
rect 3234 292544 3240 292596
rect 3292 292584 3298 292596
rect 11698 292584 11704 292596
rect 3292 292556 11704 292584
rect 3292 292544 3298 292556
rect 11698 292544 11704 292556
rect 11756 292544 11762 292596
rect 59538 289688 59544 289740
rect 59596 289728 59602 289740
rect 61194 289728 61200 289740
rect 59596 289700 61200 289728
rect 59596 289688 59602 289700
rect 61194 289688 61200 289700
rect 61252 289688 61258 289740
rect 65702 285676 65708 285728
rect 65760 285716 65766 285728
rect 68278 285716 68284 285728
rect 65760 285688 68284 285716
rect 65760 285676 65766 285688
rect 68278 285676 68284 285688
rect 68336 285676 68342 285728
rect 45738 284316 45744 284368
rect 45796 284356 45802 284368
rect 54478 284356 54484 284368
rect 45796 284328 54484 284356
rect 45796 284316 45802 284328
rect 54478 284316 54484 284328
rect 54536 284316 54542 284368
rect 57330 284316 57336 284368
rect 57388 284356 57394 284368
rect 59538 284356 59544 284368
rect 57388 284328 59544 284356
rect 57388 284316 57394 284328
rect 59538 284316 59544 284328
rect 59596 284316 59602 284368
rect 57974 282888 57980 282940
rect 58032 282928 58038 282940
rect 59998 282928 60004 282940
rect 58032 282900 60004 282928
rect 58032 282888 58038 282900
rect 59998 282888 60004 282900
rect 60056 282888 60062 282940
rect 53098 280780 53104 280832
rect 53156 280820 53162 280832
rect 57330 280820 57336 280832
rect 53156 280792 57336 280820
rect 53156 280780 53162 280792
rect 57330 280780 57336 280792
rect 57388 280780 57394 280832
rect 53834 278740 53840 278792
rect 53892 278780 53898 278792
rect 57882 278780 57888 278792
rect 53892 278752 57888 278780
rect 53892 278740 53898 278752
rect 57882 278740 57888 278752
rect 57940 278740 57946 278792
rect 61378 277380 61384 277432
rect 61436 277420 61442 277432
rect 65702 277420 65708 277432
rect 61436 277392 65708 277420
rect 61436 277380 61442 277392
rect 65702 277380 65708 277392
rect 65760 277380 65766 277432
rect 51718 276020 51724 276072
rect 51776 276060 51782 276072
rect 53098 276060 53104 276072
rect 51776 276032 53104 276060
rect 51776 276020 51782 276032
rect 53098 276020 53104 276032
rect 53156 276020 53162 276072
rect 504358 271872 504364 271924
rect 504416 271912 504422 271924
rect 579982 271912 579988 271924
rect 504416 271884 579988 271912
rect 504416 271872 504422 271884
rect 579982 271872 579988 271884
rect 580040 271872 580046 271924
rect 47578 271124 47584 271176
rect 47636 271164 47642 271176
rect 53834 271164 53840 271176
rect 47636 271136 53840 271164
rect 47636 271124 47642 271136
rect 53834 271124 53840 271136
rect 53892 271124 53898 271176
rect 3142 266364 3148 266416
rect 3200 266404 3206 266416
rect 17218 266404 17224 266416
rect 3200 266376 17224 266404
rect 3200 266364 3206 266376
rect 17218 266364 17224 266376
rect 17276 266364 17282 266416
rect 45646 263576 45652 263628
rect 45704 263616 45710 263628
rect 47578 263616 47584 263628
rect 45704 263588 47584 263616
rect 45704 263576 45710 263588
rect 47578 263576 47584 263588
rect 47636 263576 47642 263628
rect 45186 261468 45192 261520
rect 45244 261508 45250 261520
rect 61378 261508 61384 261520
rect 45244 261480 61384 261508
rect 45244 261468 45250 261480
rect 61378 261468 61384 261480
rect 61436 261468 61442 261520
rect 406378 258068 406384 258120
rect 406436 258108 406442 258120
rect 579982 258108 579988 258120
rect 406436 258080 579988 258108
rect 406436 258068 406442 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 3234 253920 3240 253972
rect 3292 253960 3298 253972
rect 25498 253960 25504 253972
rect 3292 253932 25504 253960
rect 3292 253920 3298 253932
rect 25498 253920 25504 253932
rect 25556 253920 25562 253972
rect 48222 253172 48228 253224
rect 48280 253212 48286 253224
rect 51718 253212 51724 253224
rect 48280 253184 51724 253212
rect 48280 253172 48286 253184
rect 51718 253172 51724 253184
rect 51776 253172 51782 253224
rect 45554 249432 45560 249484
rect 45612 249472 45618 249484
rect 48222 249472 48228 249484
rect 45612 249444 48228 249472
rect 45612 249432 45618 249444
rect 48222 249432 48228 249444
rect 48280 249432 48286 249484
rect 397086 244264 397092 244316
rect 397144 244304 397150 244316
rect 579982 244304 579988 244316
rect 397144 244276 579988 244304
rect 397144 244264 397150 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 45462 241340 45468 241392
rect 45520 241380 45526 241392
rect 45830 241380 45836 241392
rect 45520 241352 45836 241380
rect 45520 241340 45526 241352
rect 45830 241340 45836 241352
rect 45888 241340 45894 241392
rect 44910 240864 44916 240916
rect 44968 240904 44974 240916
rect 71774 240904 71780 240916
rect 44968 240876 71780 240904
rect 44968 240864 44974 240876
rect 71774 240864 71780 240876
rect 71832 240864 71838 240916
rect 45002 240796 45008 240848
rect 45060 240836 45066 240848
rect 88334 240836 88340 240848
rect 45060 240808 88340 240836
rect 45060 240796 45066 240808
rect 88334 240796 88340 240808
rect 88392 240796 88398 240848
rect 45094 240728 45100 240780
rect 45152 240768 45158 240780
rect 104894 240768 104900 240780
rect 45152 240740 104900 240768
rect 45152 240728 45158 240740
rect 104894 240728 104900 240740
rect 104952 240728 104958 240780
rect 3234 240116 3240 240168
rect 3292 240156 3298 240168
rect 44818 240156 44824 240168
rect 3292 240128 44824 240156
rect 3292 240116 3298 240128
rect 44818 240116 44824 240128
rect 44876 240116 44882 240168
rect 45462 239708 45468 239760
rect 45520 239748 45526 239760
rect 45922 239748 45928 239760
rect 45520 239720 45928 239748
rect 45520 239708 45526 239720
rect 45922 239708 45928 239720
rect 45980 239708 45986 239760
rect 45370 238756 45376 238808
rect 45428 238796 45434 238808
rect 45738 238796 45744 238808
rect 45428 238768 45744 238796
rect 45428 238756 45434 238768
rect 45738 238756 45744 238768
rect 45796 238756 45802 238808
rect 45830 233112 45836 233164
rect 45888 233152 45894 233164
rect 45888 233124 103514 233152
rect 45888 233112 45894 233124
rect 45646 232908 45652 232960
rect 45704 232948 45710 232960
rect 73798 232948 73804 232960
rect 45704 232920 73804 232948
rect 45704 232908 45710 232920
rect 73798 232908 73804 232920
rect 73856 232908 73862 232960
rect 103486 232404 103514 233124
rect 116394 232404 116400 232416
rect 103486 232376 116400 232404
rect 116394 232364 116400 232376
rect 116452 232364 116458 232416
rect 394786 232228 394792 232280
rect 394844 232268 394850 232280
rect 396534 232268 396540 232280
rect 394844 232240 396540 232268
rect 394844 232228 394850 232240
rect 396534 232228 396540 232240
rect 396592 232228 396598 232280
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 579798 231860 579804 231872
rect 394016 231832 579804 231860
rect 394016 231820 394022 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 45370 231072 45376 231124
rect 45428 231112 45434 231124
rect 50982 231112 50988 231124
rect 45428 231084 50988 231112
rect 45428 231072 45434 231084
rect 50982 231072 50988 231084
rect 51040 231072 51046 231124
rect 118602 231072 118608 231124
rect 118660 231112 118666 231124
rect 397638 231112 397644 231124
rect 118660 231084 397644 231112
rect 118660 231072 118666 231084
rect 397638 231072 397644 231084
rect 397696 231072 397702 231124
rect 45186 230460 45192 230512
rect 45244 230500 45250 230512
rect 46934 230500 46940 230512
rect 45244 230472 46940 230500
rect 45244 230460 45250 230472
rect 46934 230460 46940 230472
rect 46992 230460 46998 230512
rect 391934 230460 391940 230512
rect 391992 230500 391998 230512
rect 394786 230500 394792 230512
rect 391992 230472 394792 230500
rect 391992 230460 391998 230472
rect 394786 230460 394792 230472
rect 394844 230460 394850 230512
rect 174538 229848 174544 229900
rect 174596 229888 174602 229900
rect 176654 229888 176660 229900
rect 174596 229860 176660 229888
rect 174596 229848 174602 229860
rect 176654 229848 176660 229860
rect 176712 229848 176718 229900
rect 235258 228488 235264 228540
rect 235316 228528 235322 228540
rect 266538 228528 266544 228540
rect 235316 228500 266544 228528
rect 235316 228488 235322 228500
rect 266538 228488 266544 228500
rect 266596 228488 266602 228540
rect 166258 228420 166264 228472
rect 166316 228460 166322 228472
rect 296714 228460 296720 228472
rect 166316 228432 296720 228460
rect 166316 228420 166322 228432
rect 296714 228420 296720 228432
rect 296772 228420 296778 228472
rect 300118 228420 300124 228472
rect 300176 228460 300182 228472
rect 356514 228460 356520 228472
rect 300176 228432 356520 228460
rect 300176 228420 300182 228432
rect 356514 228420 356520 228432
rect 356572 228420 356578 228472
rect 50982 228352 50988 228404
rect 51040 228392 51046 228404
rect 58618 228392 58624 228404
rect 51040 228364 58624 228392
rect 51040 228352 51046 228364
rect 58618 228352 58624 228364
rect 58676 228352 58682 228404
rect 180058 228352 180064 228404
rect 180116 228392 180122 228404
rect 580166 228392 580172 228404
rect 180116 228364 580172 228392
rect 180116 228352 180122 228364
rect 580166 228352 580172 228364
rect 580224 228352 580230 228404
rect 3234 227740 3240 227792
rect 3292 227780 3298 227792
rect 40678 227780 40684 227792
rect 3292 227752 40684 227780
rect 3292 227740 3298 227752
rect 40678 227740 40684 227752
rect 40736 227740 40742 227792
rect 116394 227740 116400 227792
rect 116452 227780 116458 227792
rect 122098 227780 122104 227792
rect 116452 227752 122104 227780
rect 116452 227740 116458 227752
rect 122098 227740 122104 227752
rect 122156 227740 122162 227792
rect 233878 227740 233884 227792
rect 233936 227780 233942 227792
rect 236546 227780 236552 227792
rect 233936 227752 236552 227780
rect 233936 227740 233942 227752
rect 236546 227740 236552 227752
rect 236604 227740 236610 227792
rect 46934 227468 46940 227520
rect 46992 227508 46998 227520
rect 50338 227508 50344 227520
rect 46992 227480 50344 227508
rect 46992 227468 46998 227480
rect 50338 227468 50344 227480
rect 50396 227468 50402 227520
rect 180150 226992 180156 227044
rect 180208 227032 180214 227044
rect 580718 227032 580724 227044
rect 180208 227004 580724 227032
rect 180208 226992 180214 227004
rect 580718 226992 580724 227004
rect 580776 226992 580782 227044
rect 45646 224204 45652 224256
rect 45704 224244 45710 224256
rect 48958 224244 48964 224256
rect 45704 224216 48964 224244
rect 45704 224204 45710 224216
rect 48958 224204 48964 224216
rect 49016 224204 49022 224256
rect 73798 224204 73804 224256
rect 73856 224244 73862 224256
rect 77938 224244 77944 224256
rect 73856 224216 77944 224244
rect 73856 224204 73862 224216
rect 77938 224204 77944 224216
rect 77996 224204 78002 224256
rect 389818 223524 389824 223576
rect 389876 223564 389882 223576
rect 391934 223564 391940 223576
rect 389876 223536 391940 223564
rect 389876 223524 389882 223536
rect 391934 223524 391940 223536
rect 391992 223524 391998 223576
rect 58618 219852 58624 219904
rect 58676 219892 58682 219904
rect 64874 219892 64880 219904
rect 58676 219864 64880 219892
rect 58676 219852 58682 219864
rect 64874 219852 64880 219864
rect 64932 219852 64938 219904
rect 387794 218084 387800 218136
rect 387852 218124 387858 218136
rect 389818 218124 389824 218136
rect 387852 218096 389824 218124
rect 387852 218084 387858 218096
rect 389818 218084 389824 218096
rect 389876 218084 389882 218136
rect 48958 218016 48964 218068
rect 49016 218056 49022 218068
rect 49016 218028 49740 218056
rect 49016 218016 49022 218028
rect 49712 217988 49740 218028
rect 211798 218016 211804 218068
rect 211856 218056 211862 218068
rect 580166 218056 580172 218068
rect 211856 218028 580172 218056
rect 211856 218016 211862 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 51718 217988 51724 218000
rect 49712 217960 51724 217988
rect 51718 217948 51724 217960
rect 51776 217948 51782 218000
rect 50338 216044 50344 216096
rect 50396 216084 50402 216096
rect 65518 216084 65524 216096
rect 50396 216056 65524 216084
rect 50396 216044 50402 216056
rect 65518 216044 65524 216056
rect 65576 216044 65582 216096
rect 40678 215908 40684 215960
rect 40736 215948 40742 215960
rect 164234 215948 164240 215960
rect 40736 215920 164240 215948
rect 40736 215908 40742 215920
rect 164234 215908 164240 215920
rect 164292 215908 164298 215960
rect 64874 215296 64880 215348
rect 64932 215336 64938 215348
rect 68278 215336 68284 215348
rect 64932 215308 68284 215336
rect 64932 215296 64938 215308
rect 68278 215296 68284 215308
rect 68336 215296 68342 215348
rect 77938 215228 77944 215280
rect 77996 215268 78002 215280
rect 86218 215268 86224 215280
rect 77996 215240 86224 215268
rect 77996 215228 78002 215240
rect 86218 215228 86224 215240
rect 86276 215228 86282 215280
rect 122098 214548 122104 214600
rect 122156 214588 122162 214600
rect 135898 214588 135904 214600
rect 122156 214560 135904 214588
rect 122156 214548 122162 214560
rect 135898 214548 135904 214560
rect 135956 214548 135962 214600
rect 378318 214548 378324 214600
rect 378376 214588 378382 214600
rect 387794 214588 387800 214600
rect 378376 214560 387800 214588
rect 378376 214548 378382 214560
rect 387794 214548 387800 214560
rect 387852 214548 387858 214600
rect 3234 213936 3240 213988
rect 3292 213976 3298 213988
rect 90358 213976 90364 213988
rect 3292 213948 90364 213976
rect 3292 213936 3298 213948
rect 90358 213936 90364 213948
rect 90416 213936 90422 213988
rect 378318 212548 378324 212560
rect 376772 212520 378324 212548
rect 374914 212440 374920 212492
rect 374972 212480 374978 212492
rect 376772 212480 376800 212520
rect 378318 212508 378324 212520
rect 378376 212508 378382 212560
rect 374972 212452 376800 212480
rect 374972 212440 374978 212452
rect 370498 209788 370504 209840
rect 370556 209828 370562 209840
rect 374914 209828 374920 209840
rect 370556 209800 374920 209828
rect 370556 209788 370562 209800
rect 374914 209788 374920 209800
rect 374972 209788 374978 209840
rect 68278 207612 68284 207664
rect 68336 207652 68342 207664
rect 88242 207652 88248 207664
rect 68336 207624 88248 207652
rect 68336 207612 68342 207624
rect 88242 207612 88248 207624
rect 88300 207612 88306 207664
rect 118694 205640 118700 205692
rect 118752 205680 118758 205692
rect 580166 205680 580172 205692
rect 118752 205652 580172 205680
rect 118752 205640 118758 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 88242 203532 88248 203584
rect 88300 203572 88306 203584
rect 112438 203572 112444 203584
rect 88300 203544 112444 203572
rect 88300 203532 88306 203544
rect 112438 203532 112444 203544
rect 112496 203532 112502 203584
rect 154850 202104 154856 202156
rect 154908 202144 154914 202156
rect 235258 202144 235264 202156
rect 154908 202116 235264 202144
rect 154908 202104 154914 202116
rect 235258 202104 235264 202116
rect 235316 202104 235322 202156
rect 153194 200744 153200 200796
rect 153252 200784 153258 200796
rect 233878 200784 233884 200796
rect 153252 200756 233884 200784
rect 153252 200744 153258 200756
rect 233878 200744 233884 200756
rect 233936 200744 233942 200796
rect 148962 199384 148968 199436
rect 149020 199424 149026 199436
rect 207014 199424 207020 199436
rect 149020 199396 207020 199424
rect 149020 199384 149026 199396
rect 207014 199384 207020 199396
rect 207072 199384 207078 199436
rect 86218 199180 86224 199232
rect 86276 199220 86282 199232
rect 88794 199220 88800 199232
rect 86276 199192 88800 199220
rect 86276 199180 86282 199192
rect 88794 199180 88800 199192
rect 88852 199180 88858 199232
rect 112438 198908 112444 198960
rect 112496 198948 112502 198960
rect 115198 198948 115204 198960
rect 112496 198920 115204 198948
rect 112496 198908 112502 198920
rect 115198 198908 115204 198920
rect 115256 198908 115262 198960
rect 158898 197956 158904 198008
rect 158956 197996 158962 198008
rect 386414 197996 386420 198008
rect 158956 197968 386420 197996
rect 158956 197956 158962 197968
rect 386414 197956 386420 197968
rect 386472 197956 386478 198008
rect 151078 197412 151084 197464
rect 151136 197452 151142 197464
rect 153194 197452 153200 197464
rect 151136 197424 153200 197452
rect 151136 197412 151142 197424
rect 153194 197412 153200 197424
rect 153252 197412 153258 197464
rect 152734 197344 152740 197396
rect 152792 197384 152798 197396
rect 154850 197384 154856 197396
rect 152792 197356 154856 197384
rect 152792 197344 152798 197356
rect 154850 197344 154856 197356
rect 154908 197344 154914 197396
rect 367738 197344 367744 197396
rect 367796 197384 367802 197396
rect 370498 197384 370504 197396
rect 367796 197356 370504 197384
rect 367796 197344 367802 197356
rect 370498 197344 370504 197356
rect 370556 197344 370562 197396
rect 154482 196732 154488 196784
rect 154540 196772 154546 196784
rect 166258 196772 166264 196784
rect 154540 196744 166264 196772
rect 154540 196732 154546 196744
rect 166258 196732 166264 196744
rect 166316 196732 166322 196784
rect 147950 196664 147956 196716
rect 148008 196704 148014 196716
rect 174538 196704 174544 196716
rect 148008 196676 174544 196704
rect 148008 196664 148014 196676
rect 174538 196664 174544 196676
rect 174596 196664 174602 196716
rect 156138 196596 156144 196648
rect 156196 196636 156202 196648
rect 327074 196636 327080 196648
rect 156196 196608 327080 196636
rect 156196 196596 156202 196608
rect 327074 196596 327080 196608
rect 327132 196596 327138 196648
rect 135898 196256 135904 196308
rect 135956 196296 135962 196308
rect 138474 196296 138480 196308
rect 135956 196268 138480 196296
rect 135956 196256 135962 196268
rect 138474 196256 138480 196268
rect 138532 196256 138538 196308
rect 56594 195916 56600 195968
rect 56652 195956 56658 195968
rect 138106 195956 138112 195968
rect 56652 195928 138112 195956
rect 56652 195916 56658 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 157518 195916 157524 195968
rect 157576 195956 157582 195968
rect 300118 195956 300124 195968
rect 157576 195928 300124 195956
rect 157576 195916 157582 195928
rect 300118 195916 300124 195928
rect 300176 195916 300182 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 51718 195644 51724 195696
rect 51776 195684 51782 195696
rect 53466 195684 53472 195696
rect 51776 195656 53472 195684
rect 51776 195644 51782 195656
rect 53466 195644 53472 195656
rect 53524 195644 53530 195696
rect 115934 194556 115940 194608
rect 115992 194596 115998 194608
rect 140774 194596 140780 194608
rect 115992 194568 140780 194596
rect 115992 194556 115998 194568
rect 140774 194556 140780 194568
rect 140832 194556 140838 194608
rect 88794 194488 88800 194540
rect 88852 194528 88858 194540
rect 91738 194528 91744 194540
rect 88852 194500 91744 194528
rect 88852 194488 88858 194500
rect 91738 194488 91744 194500
rect 91796 194488 91802 194540
rect 180242 191836 180248 191888
rect 180300 191876 180306 191888
rect 579798 191876 579804 191888
rect 180300 191848 579804 191876
rect 180300 191836 180306 191848
rect 579798 191836 579804 191848
rect 579856 191836 579862 191888
rect 140774 190952 140780 191004
rect 140832 190952 140838 191004
rect 53466 190544 53472 190596
rect 53524 190584 53530 190596
rect 55858 190584 55864 190596
rect 53524 190556 55864 190584
rect 53524 190544 53530 190556
rect 55858 190544 55864 190556
rect 55916 190544 55922 190596
rect 140792 190528 140820 190952
rect 140774 190476 140780 190528
rect 140832 190476 140838 190528
rect 144730 190476 144736 190528
rect 144788 190516 144794 190528
rect 149606 190516 149612 190528
rect 144788 190488 149612 190516
rect 144788 190476 144794 190488
rect 149606 190476 149612 190488
rect 149664 190476 149670 190528
rect 140682 190408 140688 190460
rect 140740 190448 140746 190460
rect 140740 190420 140820 190448
rect 140740 190408 140746 190420
rect 140792 190256 140820 190420
rect 165430 190340 165436 190392
rect 165488 190340 165494 190392
rect 140774 190204 140780 190256
rect 140832 190204 140838 190256
rect 165448 189100 165476 190340
rect 165430 189048 165436 189100
rect 165488 189048 165494 189100
rect 3142 187688 3148 187740
rect 3200 187728 3206 187740
rect 119338 187728 119344 187740
rect 3200 187700 119344 187728
rect 3200 187688 3206 187700
rect 119338 187688 119344 187700
rect 119396 187688 119402 187740
rect 144454 180956 144460 181008
rect 144512 180996 144518 181008
rect 146018 180996 146024 181008
rect 144512 180968 146024 180996
rect 144512 180956 144518 180968
rect 146018 180956 146024 180968
rect 146076 180956 146082 181008
rect 91738 180820 91744 180872
rect 91796 180860 91802 180872
rect 95878 180860 95884 180872
rect 91796 180832 95884 180860
rect 91796 180820 91802 180832
rect 95878 180820 95884 180832
rect 95936 180820 95942 180872
rect 121454 180072 121460 180124
rect 121512 180112 121518 180124
rect 136358 180112 136364 180124
rect 121512 180084 136364 180112
rect 121512 180072 121518 180084
rect 136358 180072 136364 180084
rect 136416 180072 136422 180124
rect 135990 178848 135996 178900
rect 136048 178888 136054 178900
rect 136542 178888 136548 178900
rect 136048 178860 136548 178888
rect 136048 178848 136054 178860
rect 136542 178848 136548 178860
rect 136600 178848 136606 178900
rect 122834 178644 122840 178696
rect 122892 178684 122898 178696
rect 136450 178684 136456 178696
rect 122892 178656 136456 178684
rect 122892 178644 122898 178656
rect 136450 178644 136456 178656
rect 136508 178644 136514 178696
rect 211890 178032 211896 178084
rect 211948 178072 211954 178084
rect 579982 178072 579988 178084
rect 211948 178044 579988 178072
rect 211948 178032 211954 178044
rect 579982 178032 579988 178044
rect 580040 178032 580046 178084
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 135990 177324 135996 177336
rect 124272 177296 135996 177324
rect 124272 177284 124278 177296
rect 135990 177284 135996 177296
rect 136048 177284 136054 177336
rect 65518 177216 65524 177268
rect 65576 177256 65582 177268
rect 72418 177256 72424 177268
rect 65576 177228 72424 177256
rect 65576 177216 65582 177228
rect 72418 177216 72424 177228
rect 72476 177216 72482 177268
rect 366358 176672 366364 176724
rect 366416 176712 366422 176724
rect 367738 176712 367744 176724
rect 366416 176684 367744 176712
rect 366416 176672 366422 176684
rect 367738 176672 367744 176684
rect 367796 176672 367802 176724
rect 126974 176060 126980 176112
rect 127032 176100 127038 176112
rect 136266 176100 136272 176112
rect 127032 176072 136272 176100
rect 127032 176060 127038 176072
rect 136266 176060 136272 176072
rect 136324 176060 136330 176112
rect 149330 176032 149336 176044
rect 142126 176004 149336 176032
rect 125594 175924 125600 175976
rect 125652 175964 125658 175976
rect 136174 175964 136180 175976
rect 125652 175936 136180 175964
rect 125652 175924 125658 175936
rect 136174 175924 136180 175936
rect 136232 175924 136238 175976
rect 141602 175924 141608 175976
rect 141660 175964 141666 175976
rect 142126 175964 142154 176004
rect 149330 175992 149336 176004
rect 149388 175992 149394 176044
rect 162486 175964 162492 175976
rect 141660 175936 142154 175964
rect 154408 175936 162492 175964
rect 141660 175924 141666 175936
rect 144454 175516 144460 175568
rect 144512 175556 144518 175568
rect 149974 175556 149980 175568
rect 144512 175528 149980 175556
rect 144512 175516 144518 175528
rect 149974 175516 149980 175528
rect 150032 175516 150038 175568
rect 154408 175432 154436 175936
rect 162486 175924 162492 175936
rect 162544 175924 162550 175976
rect 154390 175380 154396 175432
rect 154448 175380 154454 175432
rect 128354 175176 128360 175228
rect 128412 175216 128418 175228
rect 136358 175216 136364 175228
rect 128412 175188 136364 175216
rect 128412 175176 128418 175188
rect 136358 175176 136364 175188
rect 136416 175176 136422 175228
rect 142062 174808 142068 174820
rect 141620 174780 142068 174808
rect 141620 174468 141648 174780
rect 142062 174768 142068 174780
rect 142120 174768 142126 174820
rect 141694 174700 141700 174752
rect 141752 174700 141758 174752
rect 144086 174700 144092 174752
rect 144144 174740 144150 174752
rect 145466 174740 145472 174752
rect 144144 174712 145472 174740
rect 144144 174700 144150 174712
rect 145466 174700 145472 174712
rect 145524 174700 145530 174752
rect 141712 174536 141740 174700
rect 152458 174632 152464 174684
rect 152516 174672 152522 174684
rect 156506 174672 156512 174684
rect 152516 174644 156512 174672
rect 152516 174632 152522 174644
rect 156506 174632 156512 174644
rect 156564 174632 156570 174684
rect 161474 174536 161480 174548
rect 141712 174508 161480 174536
rect 161474 174496 161480 174508
rect 161532 174496 161538 174548
rect 141620 174440 142154 174468
rect 142126 174332 142154 174440
rect 166994 174332 167000 174344
rect 142126 174304 167000 174332
rect 166994 174292 167000 174304
rect 167052 174292 167058 174344
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 137370 173924 137376 173936
rect 133932 173896 137376 173924
rect 133932 173884 133938 173896
rect 137370 173884 137376 173896
rect 137428 173884 137434 173936
rect 149330 172932 149336 172984
rect 149388 172972 149394 172984
rect 151446 172972 151452 172984
rect 149388 172944 151452 172972
rect 149388 172932 149394 172944
rect 151446 172932 151452 172944
rect 151504 172932 151510 172984
rect 158438 172932 158444 172984
rect 158496 172972 158502 172984
rect 159634 172972 159640 172984
rect 158496 172944 159640 172972
rect 158496 172932 158502 172944
rect 159634 172932 159640 172944
rect 159692 172932 159698 172984
rect 162486 172932 162492 172984
rect 162544 172972 162550 172984
rect 165522 172972 165528 172984
rect 162544 172944 165528 172972
rect 162544 172932 162550 172944
rect 165522 172932 165528 172944
rect 165580 172932 165586 172984
rect 131114 172524 131120 172576
rect 131172 172564 131178 172576
rect 136634 172564 136640 172576
rect 131172 172536 136640 172564
rect 131172 172524 131178 172536
rect 136634 172524 136640 172536
rect 136692 172524 136698 172576
rect 138014 172116 138020 172168
rect 138072 172156 138078 172168
rect 140774 172156 140780 172168
rect 138072 172128 140780 172156
rect 138072 172116 138078 172128
rect 140774 172116 140780 172128
rect 140832 172116 140838 172168
rect 135254 171640 135260 171692
rect 135312 171680 135318 171692
rect 138658 171680 138664 171692
rect 135312 171652 138664 171680
rect 135312 171640 135318 171652
rect 138658 171640 138664 171652
rect 138716 171640 138722 171692
rect 132494 171096 132500 171148
rect 132552 171136 132558 171148
rect 136726 171136 136732 171148
rect 132552 171108 136732 171136
rect 132552 171096 132558 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 55858 169736 55864 169788
rect 55916 169776 55922 169788
rect 55916 169748 56640 169776
rect 55916 169736 55922 169748
rect 56612 169708 56640 169748
rect 60734 169708 60740 169720
rect 56612 169680 60740 169708
rect 60734 169668 60740 169680
rect 60792 169668 60798 169720
rect 142430 166268 142436 166320
rect 142488 166308 142494 166320
rect 142614 166308 142620 166320
rect 142488 166280 142620 166308
rect 142488 166268 142494 166280
rect 142614 166268 142620 166280
rect 142672 166268 142678 166320
rect 146478 166268 146484 166320
rect 146536 166308 146542 166320
rect 147582 166308 147588 166320
rect 146536 166280 147588 166308
rect 146536 166268 146542 166280
rect 147582 166268 147588 166280
rect 147640 166268 147646 166320
rect 118510 165588 118516 165640
rect 118568 165628 118574 165640
rect 580166 165628 580172 165640
rect 118568 165600 580172 165628
rect 118568 165588 118574 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 60734 163276 60740 163328
rect 60792 163316 60798 163328
rect 66254 163316 66260 163328
rect 60792 163288 66260 163316
rect 60792 163276 60798 163288
rect 66254 163276 66260 163288
rect 66312 163276 66318 163328
rect 3142 162868 3148 162920
rect 3200 162908 3206 162920
rect 86218 162908 86224 162920
rect 3200 162880 86224 162908
rect 3200 162868 3206 162880
rect 86218 162868 86224 162880
rect 86276 162868 86282 162920
rect 72418 156612 72424 156664
rect 72476 156652 72482 156664
rect 79318 156652 79324 156664
rect 72476 156624 79324 156652
rect 72476 156612 72482 156624
rect 79318 156612 79324 156624
rect 79376 156612 79382 156664
rect 66254 155864 66260 155916
rect 66312 155904 66318 155916
rect 67634 155904 67640 155916
rect 66312 155876 67640 155904
rect 66312 155864 66318 155876
rect 67634 155864 67640 155876
rect 67692 155864 67698 155916
rect 67634 153144 67640 153196
rect 67692 153184 67698 153196
rect 72418 153184 72424 153196
rect 67692 153156 72424 153184
rect 67692 153144 67698 153156
rect 72418 153144 72424 153156
rect 72476 153144 72482 153196
rect 345658 151784 345664 151836
rect 345716 151824 345722 151836
rect 580166 151824 580172 151836
rect 345716 151796 580172 151824
rect 345716 151784 345722 151796
rect 580166 151784 580172 151796
rect 580224 151784 580230 151836
rect 79318 149676 79324 149728
rect 79376 149716 79382 149728
rect 87598 149716 87604 149728
rect 79376 149688 87604 149716
rect 79376 149676 79382 149688
rect 87598 149676 87604 149688
rect 87656 149676 87662 149728
rect 3326 149064 3332 149116
rect 3384 149104 3390 149116
rect 179414 149104 179420 149116
rect 3384 149076 179420 149104
rect 3384 149064 3390 149076
rect 179414 149064 179420 149076
rect 179472 149064 179478 149116
rect 158438 148384 158444 148436
rect 158496 148424 158502 148436
rect 164970 148424 164976 148436
rect 158496 148396 164976 148424
rect 158496 148384 158502 148396
rect 164970 148384 164976 148396
rect 165028 148384 165034 148436
rect 3050 148316 3056 148368
rect 3108 148356 3114 148368
rect 180794 148356 180800 148368
rect 3108 148328 180800 148356
rect 3108 148316 3114 148328
rect 180794 148316 180800 148328
rect 180852 148316 180858 148368
rect 25498 146888 25504 146940
rect 25556 146928 25562 146940
rect 182174 146928 182180 146940
rect 25556 146900 182180 146928
rect 25556 146888 25562 146900
rect 182174 146888 182180 146900
rect 182232 146888 182238 146940
rect 95878 146208 95884 146260
rect 95936 146248 95942 146260
rect 101398 146248 101404 146260
rect 95936 146220 101404 146248
rect 95936 146208 95942 146220
rect 101398 146208 101404 146220
rect 101456 146208 101462 146260
rect 146570 143488 146576 143540
rect 146628 143528 146634 143540
rect 148042 143528 148048 143540
rect 146628 143500 148048 143528
rect 146628 143488 146634 143500
rect 148042 143488 148048 143500
rect 148100 143488 148106 143540
rect 155218 143488 155224 143540
rect 155276 143528 155282 143540
rect 160094 143528 160100 143540
rect 155276 143500 160100 143528
rect 155276 143488 155282 143500
rect 160094 143488 160100 143500
rect 160152 143488 160158 143540
rect 165430 143488 165436 143540
rect 165488 143528 165494 143540
rect 169938 143528 169944 143540
rect 165488 143500 169944 143528
rect 165488 143488 165494 143500
rect 169938 143488 169944 143500
rect 169996 143488 170002 143540
rect 137738 143420 137744 143472
rect 137796 143460 137802 143472
rect 139578 143460 139584 143472
rect 137796 143432 139584 143460
rect 137796 143420 137802 143432
rect 139578 143420 139584 143432
rect 139636 143420 139642 143472
rect 146478 143420 146484 143472
rect 146536 143460 146542 143472
rect 149606 143460 149612 143472
rect 146536 143432 149612 143460
rect 146536 143420 146542 143432
rect 149606 143420 149612 143432
rect 149664 143420 149670 143472
rect 152458 143420 152464 143472
rect 152516 143460 152522 143472
rect 157426 143460 157432 143472
rect 152516 143432 157432 143460
rect 152516 143420 152522 143432
rect 157426 143420 157432 143432
rect 157484 143420 157490 143472
rect 164970 143420 164976 143472
rect 165028 143460 165034 143472
rect 168374 143460 168380 143472
rect 165028 143432 168380 143460
rect 165028 143420 165034 143432
rect 168374 143420 168380 143432
rect 168432 143420 168438 143472
rect 153470 143352 153476 143404
rect 153528 143392 153534 143404
rect 158990 143392 158996 143404
rect 153528 143364 158996 143392
rect 153528 143352 153534 143364
rect 158990 143352 158996 143364
rect 159048 143352 159054 143404
rect 150526 143080 150532 143132
rect 150584 143120 150590 143132
rect 154574 143120 154580 143132
rect 150584 143092 154580 143120
rect 150584 143080 150590 143092
rect 154574 143080 154580 143092
rect 154632 143080 154638 143132
rect 163590 143080 163596 143132
rect 163648 143120 163654 143132
rect 174630 143120 174636 143132
rect 163648 143092 174636 143120
rect 163648 143080 163654 143092
rect 174630 143080 174636 143092
rect 174688 143080 174694 143132
rect 144454 143012 144460 143064
rect 144512 143052 144518 143064
rect 160554 143052 160560 143064
rect 144512 143024 160560 143052
rect 144512 143012 144518 143024
rect 160554 143012 160560 143024
rect 160612 143012 160618 143064
rect 163498 143012 163504 143064
rect 163556 143052 163562 143064
rect 163556 143024 163820 143052
rect 163556 143012 163562 143024
rect 145466 142944 145472 142996
rect 145524 142984 145530 142996
rect 163682 142984 163688 142996
rect 145524 142956 163688 142984
rect 145524 142944 145530 142956
rect 163682 142944 163688 142956
rect 163740 142944 163746 142996
rect 163792 142984 163820 143024
rect 164510 143012 164516 143064
rect 164568 143052 164574 143064
rect 176194 143052 176200 143064
rect 164568 143024 176200 143052
rect 164568 143012 164574 143024
rect 176194 143012 176200 143024
rect 176252 143012 176258 143064
rect 178034 142984 178040 142996
rect 163792 142956 178040 142984
rect 178034 142944 178040 142956
rect 178092 142944 178098 142996
rect 142522 142876 142528 142928
rect 142580 142916 142586 142928
rect 173066 142916 173072 142928
rect 142580 142888 173072 142916
rect 142580 142876 142586 142888
rect 173066 142876 173072 142888
rect 173124 142876 173130 142928
rect 118326 142808 118332 142860
rect 118384 142848 118390 142860
rect 396810 142848 396816 142860
rect 118384 142820 396816 142848
rect 118384 142808 118390 142820
rect 396810 142808 396816 142820
rect 396868 142808 396874 142860
rect 142062 142196 142068 142248
rect 142120 142236 142126 142248
rect 142430 142236 142436 142248
rect 142120 142208 142436 142236
rect 142120 142196 142126 142208
rect 142430 142196 142436 142208
rect 142488 142196 142494 142248
rect 140682 142128 140688 142180
rect 140740 142168 140746 142180
rect 142246 142168 142252 142180
rect 140740 142140 142252 142168
rect 140740 142128 140746 142140
rect 142246 142128 142252 142140
rect 142304 142128 142310 142180
rect 149514 142128 149520 142180
rect 149572 142168 149578 142180
rect 152734 142168 152740 142180
rect 149572 142140 152740 142168
rect 149572 142128 149578 142140
rect 152734 142128 152740 142140
rect 152792 142128 152798 142180
rect 72418 141788 72424 141840
rect 72476 141828 72482 141840
rect 179506 141828 179512 141840
rect 72476 141800 179512 141828
rect 72476 141788 72482 141800
rect 179506 141788 179512 141800
rect 179564 141788 179570 141840
rect 117866 141720 117872 141772
rect 117924 141760 117930 141772
rect 397086 141760 397092 141772
rect 117924 141732 397092 141760
rect 117924 141720 117930 141732
rect 397086 141720 397092 141732
rect 397144 141720 397150 141772
rect 119154 141652 119160 141704
rect 119212 141692 119218 141704
rect 429194 141692 429200 141704
rect 119212 141664 429200 141692
rect 119212 141652 119218 141664
rect 429194 141652 429200 141664
rect 429252 141652 429258 141704
rect 119246 141584 119252 141636
rect 119304 141624 119310 141636
rect 494054 141624 494060 141636
rect 119304 141596 494060 141624
rect 119304 141584 119310 141596
rect 494054 141584 494060 141596
rect 494112 141584 494118 141636
rect 119062 141516 119068 141568
rect 119120 141556 119126 141568
rect 558914 141556 558920 141568
rect 119120 141528 558920 141556
rect 119120 141516 119126 141528
rect 558914 141516 558920 141528
rect 558972 141516 558978 141568
rect 118970 141448 118976 141500
rect 119028 141488 119034 141500
rect 580258 141488 580264 141500
rect 119028 141460 580264 141488
rect 119028 141448 119034 141460
rect 580258 141448 580264 141460
rect 580316 141448 580322 141500
rect 118878 141380 118884 141432
rect 118936 141420 118942 141432
rect 580350 141420 580356 141432
rect 118936 141392 580356 141420
rect 118936 141380 118942 141392
rect 580350 141380 580356 141392
rect 580408 141380 580414 141432
rect 116762 140972 116768 141024
rect 116820 141012 116826 141024
rect 182910 141012 182916 141024
rect 116820 140984 182916 141012
rect 116820 140972 116826 140984
rect 182910 140972 182916 140984
rect 182968 140972 182974 141024
rect 117130 140904 117136 140956
rect 117188 140944 117194 140956
rect 182358 140944 182364 140956
rect 117188 140916 182364 140944
rect 117188 140904 117194 140916
rect 182358 140904 182364 140916
rect 182416 140904 182422 140956
rect 116670 140836 116676 140888
rect 116728 140876 116734 140888
rect 182634 140876 182640 140888
rect 116728 140848 182640 140876
rect 116728 140836 116734 140848
rect 182634 140836 182640 140848
rect 182692 140836 182698 140888
rect 116946 140768 116952 140820
rect 117004 140808 117010 140820
rect 182450 140808 182456 140820
rect 117004 140780 182456 140808
rect 117004 140768 117010 140780
rect 182450 140768 182456 140780
rect 182508 140768 182514 140820
rect 160094 140292 160100 140344
rect 160152 140332 160158 140344
rect 180426 140332 180432 140344
rect 160152 140304 180432 140332
rect 160152 140292 160158 140304
rect 180426 140292 180432 140304
rect 180484 140292 180490 140344
rect 118142 140224 118148 140276
rect 118200 140264 118206 140276
rect 396994 140264 397000 140276
rect 118200 140236 397000 140264
rect 118200 140224 118206 140236
rect 396994 140224 397000 140236
rect 397052 140224 397058 140276
rect 117958 140156 117964 140208
rect 118016 140196 118022 140208
rect 396902 140196 396908 140208
rect 118016 140168 396908 140196
rect 118016 140156 118022 140168
rect 396902 140156 396908 140168
rect 396960 140156 396966 140208
rect 118786 140088 118792 140140
rect 118844 140128 118850 140140
rect 580626 140128 580632 140140
rect 118844 140100 580632 140128
rect 118844 140088 118850 140100
rect 580626 140088 580632 140100
rect 580684 140088 580690 140140
rect 117774 140020 117780 140072
rect 117832 140060 117838 140072
rect 580902 140060 580908 140072
rect 117832 140032 580908 140060
rect 117832 140020 117838 140032
rect 580902 140020 580908 140032
rect 580960 140020 580966 140072
rect 179506 139816 179512 139868
rect 179564 139856 179570 139868
rect 180978 139856 180984 139868
rect 179564 139828 180984 139856
rect 179564 139816 179570 139828
rect 180978 139816 180984 139828
rect 181036 139816 181042 139868
rect 120534 139748 120540 139800
rect 120592 139788 120598 139800
rect 182266 139788 182272 139800
rect 120592 139760 182272 139788
rect 120592 139748 120598 139760
rect 182266 139748 182272 139760
rect 182324 139748 182330 139800
rect 120626 139680 120632 139732
rect 120684 139720 120690 139732
rect 182818 139720 182824 139732
rect 120684 139692 182824 139720
rect 120684 139680 120690 139692
rect 182818 139680 182824 139692
rect 182876 139680 182882 139732
rect 117222 139612 117228 139664
rect 117280 139652 117286 139664
rect 183002 139652 183008 139664
rect 117280 139624 183008 139652
rect 117280 139612 117286 139624
rect 183002 139612 183008 139624
rect 183060 139612 183066 139664
rect 116394 139544 116400 139596
rect 116452 139584 116458 139596
rect 182726 139584 182732 139596
rect 116452 139556 182732 139584
rect 116452 139544 116458 139556
rect 182726 139544 182732 139556
rect 182784 139544 182790 139596
rect 116854 139476 116860 139528
rect 116912 139516 116918 139528
rect 182542 139516 182548 139528
rect 116912 139488 182548 139516
rect 116912 139476 116918 139488
rect 182542 139476 182548 139488
rect 182600 139476 182606 139528
rect 3234 139408 3240 139460
rect 3292 139448 3298 139460
rect 179506 139448 179512 139460
rect 3292 139420 179512 139448
rect 3292 139408 3298 139420
rect 179506 139408 179512 139420
rect 179564 139408 179570 139460
rect 361574 138048 361580 138100
rect 361632 138088 361638 138100
rect 366358 138088 366364 138100
rect 361632 138060 366364 138088
rect 361632 138048 361638 138060
rect 366358 138048 366364 138060
rect 366416 138048 366422 138100
rect 189718 137980 189724 138032
rect 189776 138020 189782 138032
rect 580166 138020 580172 138032
rect 189776 137992 580172 138020
rect 189776 137980 189782 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 101398 137232 101404 137284
rect 101456 137272 101462 137284
rect 106918 137272 106924 137284
rect 101456 137244 106924 137272
rect 101456 137232 101462 137244
rect 106918 137232 106924 137244
rect 106976 137232 106982 137284
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 116578 136660 116584 136672
rect 3384 136632 116584 136660
rect 3384 136620 3390 136632
rect 116578 136620 116584 136632
rect 116636 136620 116642 136672
rect 3142 136552 3148 136604
rect 3200 136592 3206 136604
rect 117222 136592 117228 136604
rect 3200 136564 117228 136592
rect 3200 136552 3206 136564
rect 117222 136552 117228 136564
rect 117280 136592 117286 136604
rect 118418 136592 118424 136604
rect 117280 136564 118424 136592
rect 117280 136552 117286 136564
rect 118418 136552 118424 136564
rect 118476 136552 118482 136604
rect 23474 136484 23480 136536
rect 23532 136524 23538 136536
rect 118234 136524 118240 136536
rect 23532 136496 118240 136524
rect 23532 136484 23538 136496
rect 118234 136484 118240 136496
rect 118292 136484 118298 136536
rect 360838 135260 360844 135312
rect 360896 135300 360902 135312
rect 361574 135300 361580 135312
rect 360896 135272 361580 135300
rect 360896 135260 360902 135272
rect 361574 135260 361580 135272
rect 361632 135260 361638 135312
rect 18598 135192 18604 135244
rect 18656 135232 18662 135244
rect 118418 135232 118424 135244
rect 18656 135204 118424 135232
rect 18656 135192 18662 135204
rect 118418 135192 118424 135204
rect 118476 135192 118482 135244
rect 117866 134852 117872 134904
rect 117924 134892 117930 134904
rect 118418 134892 118424 134904
rect 117924 134864 118424 134892
rect 117924 134852 117930 134864
rect 118418 134852 118424 134864
rect 118476 134852 118482 134904
rect 21358 133832 21364 133884
rect 21416 133872 21422 133884
rect 117130 133872 117136 133884
rect 21416 133844 117136 133872
rect 21416 133832 21422 133844
rect 117130 133832 117136 133844
rect 117188 133832 117194 133884
rect 31018 132404 31024 132456
rect 31076 132444 31082 132456
rect 116946 132444 116952 132456
rect 31076 132416 116952 132444
rect 31076 132404 31082 132416
rect 116946 132404 116952 132416
rect 117004 132404 117010 132456
rect 32398 132336 32404 132388
rect 32456 132376 32462 132388
rect 116854 132376 116860 132388
rect 32456 132348 116860 132376
rect 32456 132336 32462 132348
rect 116854 132336 116860 132348
rect 116912 132336 116918 132388
rect 359458 131112 359464 131164
rect 359516 131152 359522 131164
rect 360838 131152 360844 131164
rect 359516 131124 360844 131152
rect 359516 131112 359522 131124
rect 360838 131112 360844 131124
rect 360896 131112 360902 131164
rect 22738 131044 22744 131096
rect 22796 131084 22802 131096
rect 116670 131084 116676 131096
rect 22796 131056 116676 131084
rect 22796 131044 22802 131056
rect 116670 131044 116676 131056
rect 116728 131044 116734 131096
rect 115198 130364 115204 130416
rect 115256 130404 115262 130416
rect 120718 130404 120724 130416
rect 115256 130376 120724 130404
rect 115256 130364 115262 130376
rect 120718 130364 120724 130376
rect 120776 130364 120782 130416
rect 28258 129684 28264 129736
rect 28316 129724 28322 129736
rect 116394 129724 116400 129736
rect 28316 129696 116400 129724
rect 28316 129684 28322 129696
rect 116394 129684 116400 129696
rect 116452 129724 116458 129736
rect 117314 129724 117320 129736
rect 116452 129696 117320 129724
rect 116452 129684 116458 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 4062 128256 4068 128308
rect 4120 128296 4126 128308
rect 116762 128296 116768 128308
rect 4120 128268 116768 128296
rect 4120 128256 4126 128268
rect 116762 128256 116768 128268
rect 116820 128296 116826 128308
rect 117314 128296 117320 128308
rect 116820 128268 117320 128296
rect 116820 128256 116826 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 90358 126216 90364 126268
rect 90416 126256 90422 126268
rect 117314 126256 117320 126268
rect 90416 126228 117320 126256
rect 90416 126216 90422 126228
rect 117314 126216 117320 126228
rect 117372 126216 117378 126268
rect 180334 125604 180340 125656
rect 180392 125644 180398 125656
rect 580166 125644 580172 125656
rect 180392 125616 580172 125644
rect 180392 125604 180398 125616
rect 580166 125604 580172 125616
rect 580224 125604 580230 125656
rect 7650 123428 7656 123480
rect 7708 123468 7714 123480
rect 117774 123468 117780 123480
rect 7708 123440 117780 123468
rect 7708 123428 7714 123440
rect 117774 123428 117780 123440
rect 117832 123428 117838 123480
rect 17310 122068 17316 122120
rect 17368 122108 17374 122120
rect 117682 122108 117688 122120
rect 17368 122080 117688 122108
rect 17368 122068 17374 122080
rect 117682 122068 117688 122080
rect 117740 122068 117746 122120
rect 106918 121456 106924 121508
rect 106976 121496 106982 121508
rect 109678 121496 109684 121508
rect 106976 121468 109684 121496
rect 106976 121456 106982 121468
rect 109678 121456 109684 121468
rect 109736 121456 109742 121508
rect 86218 121388 86224 121440
rect 86276 121428 86282 121440
rect 117314 121428 117320 121440
rect 86276 121400 117320 121428
rect 86276 121388 86282 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 180426 120776 180432 120828
rect 180484 120816 180490 120828
rect 182174 120816 182180 120828
rect 180484 120788 182180 120816
rect 180484 120776 180490 120788
rect 182174 120776 182180 120788
rect 182232 120776 182238 120828
rect 6178 120096 6184 120148
rect 6236 120136 6242 120148
rect 117406 120136 117412 120148
rect 6236 120108 117412 120136
rect 6236 120096 6242 120108
rect 117406 120096 117412 120108
rect 117464 120096 117470 120148
rect 17218 118600 17224 118652
rect 17276 118640 17282 118652
rect 117314 118640 117320 118652
rect 17276 118612 117320 118640
rect 17276 118600 17282 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 87598 118532 87604 118584
rect 87656 118572 87662 118584
rect 92474 118572 92480 118584
rect 87656 118544 92480 118572
rect 87656 118532 87662 118544
rect 92474 118532 92480 118544
rect 92532 118532 92538 118584
rect 14458 117240 14464 117292
rect 14516 117280 14522 117292
rect 117406 117280 117412 117292
rect 14516 117252 117412 117280
rect 14516 117240 14522 117252
rect 117406 117240 117412 117252
rect 117464 117240 117470 117292
rect 26878 117172 26884 117224
rect 26936 117212 26942 117224
rect 117314 117212 117320 117224
rect 26936 117184 117320 117212
rect 26936 117172 26942 117184
rect 117314 117172 117320 117184
rect 117372 117172 117378 117224
rect 10318 115880 10324 115932
rect 10376 115920 10382 115932
rect 117314 115920 117320 115932
rect 10376 115892 117320 115920
rect 10376 115880 10382 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 92474 114520 92480 114572
rect 92532 114560 92538 114572
rect 95878 114560 95884 114572
rect 92532 114532 95884 114560
rect 92532 114520 92538 114532
rect 95878 114520 95884 114532
rect 95936 114520 95942 114572
rect 13078 114452 13084 114504
rect 13136 114492 13142 114504
rect 117314 114492 117320 114504
rect 13136 114464 117320 114492
rect 13136 114452 13142 114464
rect 117314 114452 117320 114464
rect 117372 114452 117378 114504
rect 8938 113092 8944 113144
rect 8996 113132 9002 113144
rect 117314 113132 117320 113144
rect 8996 113104 117320 113132
rect 8996 113092 9002 113104
rect 117314 113092 117320 113104
rect 117372 113092 117378 113144
rect 180426 111800 180432 111852
rect 180484 111840 180490 111852
rect 580166 111840 580172 111852
rect 180484 111812 580172 111840
rect 180484 111800 180490 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 4890 111732 4896 111784
rect 4948 111772 4954 111784
rect 117314 111772 117320 111784
rect 4948 111744 117320 111772
rect 4948 111732 4954 111744
rect 117314 111732 117320 111744
rect 117372 111732 117378 111784
rect 7558 111664 7564 111716
rect 7616 111704 7622 111716
rect 117406 111704 117412 111716
rect 7616 111676 117412 111704
rect 7616 111664 7622 111676
rect 117406 111664 117412 111676
rect 117464 111664 117470 111716
rect 3142 111460 3148 111512
rect 3200 111500 3206 111512
rect 6178 111500 6184 111512
rect 3200 111472 6184 111500
rect 3200 111460 3206 111472
rect 6178 111460 6184 111472
rect 6236 111460 6242 111512
rect 357434 110440 357440 110492
rect 357492 110480 357498 110492
rect 359458 110480 359464 110492
rect 357492 110452 359464 110480
rect 357492 110440 357498 110452
rect 359458 110440 359464 110452
rect 359516 110440 359522 110492
rect 4798 110372 4804 110424
rect 4856 110412 4862 110424
rect 117314 110412 117320 110424
rect 4856 110384 117320 110412
rect 4856 110372 4862 110384
rect 117314 110372 117320 110384
rect 117372 110372 117378 110424
rect 182818 109692 182824 109744
rect 182876 109732 182882 109744
rect 211798 109732 211804 109744
rect 182876 109704 211804 109732
rect 182876 109692 182882 109704
rect 211798 109692 211804 109704
rect 211856 109692 211862 109744
rect 40034 108944 40040 108996
rect 40092 108984 40098 108996
rect 117314 108984 117320 108996
rect 40092 108956 117320 108984
rect 40092 108944 40098 108956
rect 117314 108944 117320 108956
rect 117372 108944 117378 108996
rect 45094 107584 45100 107636
rect 45152 107624 45158 107636
rect 117314 107624 117320 107636
rect 45152 107596 117320 107624
rect 45152 107584 45158 107596
rect 117314 107584 117320 107596
rect 117372 107584 117378 107636
rect 183278 107584 183284 107636
rect 183336 107624 183342 107636
rect 357434 107624 357440 107636
rect 183336 107596 357440 107624
rect 183336 107584 183342 107596
rect 357434 107584 357440 107596
rect 357492 107584 357498 107636
rect 45278 106224 45284 106276
rect 45336 106264 45342 106276
rect 117314 106264 117320 106276
rect 45336 106236 117320 106264
rect 45336 106224 45342 106236
rect 117314 106224 117320 106236
rect 117372 106224 117378 106276
rect 183278 106224 183284 106276
rect 183336 106264 183342 106276
rect 396442 106264 396448 106276
rect 183336 106236 396448 106264
rect 183336 106224 183342 106236
rect 396442 106224 396448 106236
rect 396500 106224 396506 106276
rect 44634 106156 44640 106208
rect 44692 106196 44698 106208
rect 117406 106196 117412 106208
rect 44692 106168 117412 106196
rect 44692 106156 44698 106168
rect 117406 106156 117412 106168
rect 117464 106156 117470 106208
rect 44726 104796 44732 104848
rect 44784 104836 44790 104848
rect 117314 104836 117320 104848
rect 44784 104808 117320 104836
rect 44784 104796 44790 104808
rect 117314 104796 117320 104808
rect 117372 104796 117378 104848
rect 183278 104796 183284 104848
rect 183336 104836 183342 104848
rect 404998 104836 405004 104848
rect 183336 104808 405004 104836
rect 183336 104796 183342 104808
rect 404998 104796 405004 104808
rect 405056 104796 405062 104848
rect 95878 104728 95884 104780
rect 95936 104768 95942 104780
rect 99558 104768 99564 104780
rect 95936 104740 99564 104768
rect 95936 104728 95942 104740
rect 99558 104728 99564 104740
rect 99616 104728 99622 104780
rect 183278 103436 183284 103488
rect 183336 103476 183342 103488
rect 403618 103476 403624 103488
rect 183336 103448 403624 103476
rect 183336 103436 183342 103448
rect 403618 103436 403624 103448
rect 403676 103436 403682 103488
rect 183278 102076 183284 102128
rect 183336 102116 183342 102128
rect 400858 102116 400864 102128
rect 183336 102088 400864 102116
rect 183336 102076 183342 102088
rect 400858 102076 400864 102088
rect 400916 102076 400922 102128
rect 109678 101396 109684 101448
rect 109736 101436 109742 101448
rect 119430 101436 119436 101448
rect 109736 101408 119436 101436
rect 109736 101396 109742 101408
rect 119430 101396 119436 101408
rect 119488 101396 119494 101448
rect 183186 100648 183192 100700
rect 183244 100688 183250 100700
rect 399478 100688 399484 100700
rect 183244 100660 399484 100688
rect 183244 100648 183250 100660
rect 399478 100648 399484 100660
rect 399536 100648 399542 100700
rect 238018 99356 238024 99408
rect 238076 99396 238082 99408
rect 580166 99396 580172 99408
rect 238076 99368 580172 99396
rect 238076 99356 238082 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 183186 99288 183192 99340
rect 183244 99328 183250 99340
rect 417418 99328 417424 99340
rect 183244 99300 417424 99328
rect 183244 99288 183250 99300
rect 417418 99288 417424 99300
rect 417476 99288 417482 99340
rect 99558 97928 99564 97980
rect 99616 97968 99622 97980
rect 102778 97968 102784 97980
rect 99616 97940 102784 97968
rect 99616 97928 99622 97940
rect 102778 97928 102784 97940
rect 102836 97928 102842 97980
rect 183186 97928 183192 97980
rect 183244 97968 183250 97980
rect 414658 97968 414664 97980
rect 183244 97940 414664 97968
rect 183244 97928 183250 97940
rect 414658 97928 414664 97940
rect 414716 97928 414722 97980
rect 183186 96568 183192 96620
rect 183244 96608 183250 96620
rect 413278 96608 413284 96620
rect 183244 96580 413284 96608
rect 183244 96568 183250 96580
rect 413278 96568 413284 96580
rect 413336 96568 413342 96620
rect 183462 95140 183468 95192
rect 183520 95180 183526 95192
rect 522298 95180 522304 95192
rect 183520 95152 522304 95180
rect 183520 95140 183526 95152
rect 522298 95140 522304 95152
rect 522356 95140 522362 95192
rect 183462 93780 183468 93832
rect 183520 93820 183526 93832
rect 409138 93820 409144 93832
rect 183520 93792 409144 93820
rect 183520 93780 183526 93792
rect 409138 93780 409144 93792
rect 409196 93780 409202 93832
rect 183462 92420 183468 92472
rect 183520 92460 183526 92472
rect 418798 92460 418804 92472
rect 183520 92432 418804 92460
rect 183520 92420 183526 92432
rect 418798 92420 418804 92432
rect 418856 92420 418862 92472
rect 102778 90992 102784 91044
rect 102836 91032 102842 91044
rect 105630 91032 105636 91044
rect 102836 91004 105636 91032
rect 102836 90992 102842 91004
rect 105630 90992 105636 91004
rect 105688 90992 105694 91044
rect 183462 90992 183468 91044
rect 183520 91032 183526 91044
rect 407758 91032 407764 91044
rect 183520 91004 407764 91032
rect 183520 90992 183526 91004
rect 407758 90992 407764 91004
rect 407816 90992 407822 91044
rect 182266 89632 182272 89684
rect 182324 89672 182330 89684
rect 406378 89672 406384 89684
rect 182324 89644 406384 89672
rect 182324 89632 182330 89644
rect 406378 89632 406384 89644
rect 406436 89632 406442 89684
rect 182726 87592 182732 87644
rect 182784 87632 182790 87644
rect 211890 87632 211896 87644
rect 182784 87604 211896 87632
rect 182784 87592 182790 87604
rect 211890 87592 211896 87604
rect 211948 87592 211954 87644
rect 105630 86912 105636 86964
rect 105688 86952 105694 86964
rect 108114 86952 108120 86964
rect 105688 86924 108120 86952
rect 105688 86912 105694 86924
rect 108114 86912 108120 86924
rect 108172 86912 108178 86964
rect 179966 85552 179972 85604
rect 180024 85592 180030 85604
rect 580166 85592 580172 85604
rect 180024 85564 580172 85592
rect 180024 85552 180030 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 182726 85484 182732 85536
rect 182784 85524 182790 85536
rect 189718 85524 189724 85536
rect 182784 85496 189724 85524
rect 182784 85484 182790 85496
rect 189718 85484 189724 85496
rect 189776 85484 189782 85536
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 120626 84232 120632 84244
rect 3200 84204 120632 84232
rect 3200 84192 3206 84204
rect 120626 84192 120632 84204
rect 120684 84192 120690 84244
rect 182726 84124 182732 84176
rect 182784 84164 182790 84176
rect 238018 84164 238024 84176
rect 182784 84136 238024 84164
rect 182784 84124 182790 84136
rect 238018 84124 238024 84136
rect 238076 84124 238082 84176
rect 178954 81200 178960 81252
rect 179012 81240 179018 81252
rect 180334 81240 180340 81252
rect 179012 81212 180340 81240
rect 179012 81200 179018 81212
rect 180334 81200 180340 81212
rect 180392 81200 180398 81252
rect 108114 80724 108120 80776
rect 108172 80764 108178 80776
rect 120074 80764 120080 80776
rect 108172 80736 120080 80764
rect 108172 80724 108178 80736
rect 120074 80724 120080 80736
rect 120132 80724 120138 80776
rect 178954 80764 178960 80776
rect 177776 80736 178960 80764
rect 177776 80696 177804 80736
rect 178954 80724 178960 80736
rect 179012 80724 179018 80776
rect 345658 80764 345664 80776
rect 181456 80736 345664 80764
rect 178586 80696 178592 80708
rect 168346 80668 177804 80696
rect 177868 80668 178592 80696
rect 118510 80588 118516 80640
rect 118568 80628 118574 80640
rect 168346 80628 168374 80668
rect 118568 80600 168374 80628
rect 118568 80588 118574 80600
rect 118602 80520 118608 80572
rect 118660 80560 118666 80572
rect 118660 80532 168374 80560
rect 118660 80520 118666 80532
rect 168346 80492 168374 80532
rect 174446 80520 174452 80572
rect 174504 80560 174510 80572
rect 177868 80560 177896 80668
rect 178586 80656 178592 80668
rect 178644 80656 178650 80708
rect 179966 80696 179972 80708
rect 179386 80668 179972 80696
rect 179386 80628 179414 80668
rect 179966 80656 179972 80668
rect 180024 80656 180030 80708
rect 174504 80532 177896 80560
rect 178006 80600 179414 80628
rect 174504 80520 174510 80532
rect 178006 80492 178034 80600
rect 168346 80464 178034 80492
rect 174446 80424 174452 80436
rect 161446 80396 174452 80424
rect 161446 80356 161474 80396
rect 174446 80384 174452 80396
rect 174504 80384 174510 80436
rect 175274 80384 175280 80436
rect 175332 80424 175338 80436
rect 181456 80424 181484 80736
rect 345658 80724 345664 80736
rect 345716 80724 345722 80776
rect 580534 80696 580540 80708
rect 175332 80396 181484 80424
rect 186286 80668 580540 80696
rect 175332 80384 175338 80396
rect 154546 80328 161474 80356
rect 125566 80192 153194 80220
rect 11698 79976 11704 80028
rect 11756 80016 11762 80028
rect 125566 80016 125594 80192
rect 11756 79988 125594 80016
rect 126118 80124 132494 80152
rect 11756 79976 11762 79988
rect 125732 79948 125738 79960
rect 124186 79920 125738 79948
rect 3878 79840 3884 79892
rect 3936 79880 3942 79892
rect 3936 79852 123524 79880
rect 3936 79840 3942 79852
rect 3694 79704 3700 79756
rect 3752 79744 3758 79756
rect 3752 79716 120580 79744
rect 3752 79704 3758 79716
rect 3510 79568 3516 79620
rect 3568 79608 3574 79620
rect 3568 79580 120488 79608
rect 3568 79568 3574 79580
rect 116578 79092 116584 79144
rect 116636 79132 116642 79144
rect 120460 79132 120488 79580
rect 120552 79200 120580 79716
rect 123496 79336 123524 79852
rect 123662 79840 123668 79892
rect 123720 79880 123726 79892
rect 124186 79880 124214 79920
rect 125732 79908 125738 79920
rect 125790 79908 125796 79960
rect 126008 79908 126014 79960
rect 126066 79908 126072 79960
rect 123720 79852 124214 79880
rect 123720 79840 123726 79852
rect 125502 79840 125508 79892
rect 125560 79880 125566 79892
rect 125824 79880 125830 79892
rect 125560 79852 125830 79880
rect 125560 79840 125566 79852
rect 125824 79840 125830 79852
rect 125882 79840 125888 79892
rect 125042 79772 125048 79824
rect 125100 79812 125106 79824
rect 126026 79812 126054 79908
rect 125100 79784 126054 79812
rect 125100 79772 125106 79784
rect 125134 79636 125140 79688
rect 125192 79676 125198 79688
rect 126118 79676 126146 80124
rect 127314 79988 128262 80016
rect 126192 79908 126198 79960
rect 126250 79908 126256 79960
rect 126284 79908 126290 79960
rect 126342 79908 126348 79960
rect 126376 79908 126382 79960
rect 126434 79908 126440 79960
rect 126468 79908 126474 79960
rect 126526 79908 126532 79960
rect 126652 79908 126658 79960
rect 126710 79908 126716 79960
rect 126836 79908 126842 79960
rect 126894 79908 126900 79960
rect 125192 79648 126146 79676
rect 125192 79636 125198 79648
rect 125870 79568 125876 79620
rect 125928 79608 125934 79620
rect 126210 79608 126238 79908
rect 126302 79824 126330 79908
rect 126284 79772 126290 79824
rect 126342 79772 126348 79824
rect 126394 79688 126422 79908
rect 126330 79636 126336 79688
rect 126388 79648 126422 79688
rect 126388 79636 126394 79648
rect 125928 79580 126238 79608
rect 125928 79568 125934 79580
rect 125686 79432 125692 79484
rect 125744 79472 125750 79484
rect 126486 79472 126514 79908
rect 126670 79824 126698 79908
rect 126670 79784 126704 79824
rect 126698 79772 126704 79784
rect 126756 79772 126762 79824
rect 126854 79756 126882 79908
rect 127204 79880 127210 79892
rect 127176 79840 127210 79880
rect 127262 79840 127268 79892
rect 127020 79772 127026 79824
rect 127078 79812 127084 79824
rect 127078 79772 127112 79812
rect 126790 79704 126796 79756
rect 126848 79716 126882 79756
rect 126848 79704 126854 79716
rect 127084 79688 127112 79772
rect 127176 79756 127204 79840
rect 127314 79756 127342 79988
rect 128234 79960 128262 79988
rect 132466 79960 132494 80124
rect 145898 80124 150388 80152
rect 137710 80056 142154 80084
rect 132834 79988 133782 80016
rect 132834 79960 132862 79988
rect 127480 79908 127486 79960
rect 127538 79908 127544 79960
rect 127848 79908 127854 79960
rect 127906 79908 127912 79960
rect 127940 79908 127946 79960
rect 127998 79908 128004 79960
rect 128216 79908 128222 79960
rect 128274 79908 128280 79960
rect 128400 79908 128406 79960
rect 128458 79908 128464 79960
rect 128492 79908 128498 79960
rect 128550 79908 128556 79960
rect 129044 79908 129050 79960
rect 129102 79908 129108 79960
rect 129136 79908 129142 79960
rect 129194 79908 129200 79960
rect 129504 79948 129510 79960
rect 129476 79908 129510 79948
rect 129562 79908 129568 79960
rect 129596 79908 129602 79960
rect 129654 79908 129660 79960
rect 130148 79908 130154 79960
rect 130206 79908 130212 79960
rect 130240 79908 130246 79960
rect 130298 79908 130304 79960
rect 130700 79908 130706 79960
rect 130758 79908 130764 79960
rect 130884 79908 130890 79960
rect 130942 79908 130948 79960
rect 130976 79908 130982 79960
rect 131034 79908 131040 79960
rect 131068 79908 131074 79960
rect 131126 79948 131132 79960
rect 131252 79948 131258 79960
rect 131126 79908 131160 79948
rect 127388 79772 127394 79824
rect 127446 79772 127452 79824
rect 127158 79704 127164 79756
rect 127216 79704 127222 79756
rect 127250 79704 127256 79756
rect 127308 79716 127342 79756
rect 127308 79704 127314 79716
rect 127406 79688 127434 79772
rect 127498 79756 127526 79908
rect 127866 79756 127894 79908
rect 127498 79716 127532 79756
rect 127526 79704 127532 79716
rect 127584 79704 127590 79756
rect 127802 79704 127808 79756
rect 127860 79716 127894 79756
rect 127860 79704 127866 79716
rect 127066 79636 127072 79688
rect 127124 79636 127130 79688
rect 127342 79636 127348 79688
rect 127400 79648 127434 79688
rect 127958 79676 127986 79908
rect 128124 79840 128130 79892
rect 128182 79840 128188 79892
rect 128142 79756 128170 79840
rect 128418 79812 128446 79908
rect 128372 79784 128446 79812
rect 128372 79756 128400 79784
rect 128142 79716 128176 79756
rect 128170 79704 128176 79716
rect 128228 79704 128234 79756
rect 128354 79704 128360 79756
rect 128412 79704 128418 79756
rect 128510 79744 128538 79908
rect 128584 79840 128590 79892
rect 128642 79840 128648 79892
rect 128860 79840 128866 79892
rect 128918 79840 128924 79892
rect 128464 79716 128538 79744
rect 128464 79688 128492 79716
rect 128602 79688 128630 79840
rect 128768 79772 128774 79824
rect 128826 79772 128832 79824
rect 128786 79688 128814 79772
rect 127958 79648 128400 79676
rect 127400 79636 127406 79648
rect 128372 79540 128400 79648
rect 128446 79636 128452 79688
rect 128504 79636 128510 79688
rect 128538 79636 128544 79688
rect 128596 79648 128630 79688
rect 128596 79636 128602 79648
rect 128722 79636 128728 79688
rect 128780 79648 128814 79688
rect 128780 79636 128786 79648
rect 128878 79620 128906 79840
rect 128952 79772 128958 79824
rect 129010 79772 129016 79824
rect 128814 79568 128820 79620
rect 128872 79580 128906 79620
rect 128872 79568 128878 79580
rect 128970 79552 128998 79772
rect 129062 79688 129090 79908
rect 129154 79880 129182 79908
rect 129154 79852 129228 79880
rect 129200 79824 129228 79852
rect 129320 79840 129326 79892
rect 129378 79840 129384 79892
rect 129182 79772 129188 79824
rect 129240 79772 129246 79824
rect 129338 79688 129366 79840
rect 129062 79648 129096 79688
rect 129090 79636 129096 79648
rect 129148 79636 129154 79688
rect 129274 79636 129280 79688
rect 129332 79648 129366 79688
rect 129332 79636 129338 79648
rect 127774 79512 128400 79540
rect 125744 79444 126514 79472
rect 125744 79432 125750 79444
rect 127618 79432 127624 79484
rect 127676 79472 127682 79484
rect 127774 79472 127802 79512
rect 128906 79500 128912 79552
rect 128964 79512 128998 79552
rect 128964 79500 128970 79512
rect 127676 79444 127802 79472
rect 127676 79432 127682 79444
rect 128998 79432 129004 79484
rect 129056 79472 129062 79484
rect 129476 79472 129504 79908
rect 129614 79620 129642 79908
rect 129780 79840 129786 79892
rect 129838 79840 129844 79892
rect 129798 79688 129826 79840
rect 130166 79824 130194 79908
rect 129964 79772 129970 79824
rect 130022 79772 130028 79824
rect 130102 79772 130108 79824
rect 130160 79784 130194 79824
rect 130160 79772 130166 79784
rect 129734 79636 129740 79688
rect 129792 79648 129826 79688
rect 129982 79688 130010 79772
rect 129982 79648 130016 79688
rect 129792 79636 129798 79648
rect 130010 79636 130016 79648
rect 130068 79636 130074 79688
rect 129550 79568 129556 79620
rect 129608 79580 129642 79620
rect 130258 79608 130286 79908
rect 130424 79840 130430 79892
rect 130482 79840 130488 79892
rect 130608 79840 130614 79892
rect 130666 79840 130672 79892
rect 129844 79580 130286 79608
rect 129608 79568 129614 79580
rect 129844 79552 129872 79580
rect 129826 79500 129832 79552
rect 129884 79500 129890 79552
rect 129056 79444 129504 79472
rect 129056 79432 129062 79444
rect 129918 79432 129924 79484
rect 129976 79472 129982 79484
rect 130442 79472 130470 79840
rect 130626 79744 130654 79840
rect 130580 79716 130654 79744
rect 130580 79620 130608 79716
rect 130718 79688 130746 79908
rect 130792 79840 130798 79892
rect 130850 79840 130856 79892
rect 130654 79636 130660 79688
rect 130712 79648 130746 79688
rect 130712 79636 130718 79648
rect 130562 79568 130568 79620
rect 130620 79568 130626 79620
rect 129976 79444 130470 79472
rect 129976 79432 129982 79444
rect 130286 79364 130292 79416
rect 130344 79404 130350 79416
rect 130810 79404 130838 79840
rect 130902 79824 130930 79908
rect 130884 79772 130890 79824
rect 130942 79772 130948 79824
rect 130994 79688 131022 79908
rect 130930 79636 130936 79688
rect 130988 79648 131022 79688
rect 130988 79636 130994 79648
rect 131132 79620 131160 79908
rect 131224 79908 131258 79948
rect 131310 79908 131316 79960
rect 131436 79948 131442 79960
rect 131362 79920 131442 79948
rect 131224 79688 131252 79908
rect 131362 79756 131390 79920
rect 131436 79908 131442 79920
rect 131494 79908 131500 79960
rect 131528 79908 131534 79960
rect 131586 79908 131592 79960
rect 131620 79908 131626 79960
rect 131678 79908 131684 79960
rect 131804 79908 131810 79960
rect 131862 79908 131868 79960
rect 132264 79908 132270 79960
rect 132322 79908 132328 79960
rect 132356 79908 132362 79960
rect 132414 79908 132420 79960
rect 132448 79908 132454 79960
rect 132506 79908 132512 79960
rect 132816 79908 132822 79960
rect 132874 79908 132880 79960
rect 133184 79948 133190 79960
rect 133018 79920 133190 79948
rect 131546 79880 131574 79908
rect 131298 79704 131304 79756
rect 131356 79716 131390 79756
rect 131500 79852 131574 79880
rect 131356 79704 131362 79716
rect 131206 79636 131212 79688
rect 131264 79636 131270 79688
rect 131500 79620 131528 79852
rect 131638 79824 131666 79908
rect 131574 79772 131580 79824
rect 131632 79784 131666 79824
rect 131632 79772 131638 79784
rect 131114 79568 131120 79620
rect 131172 79568 131178 79620
rect 131482 79568 131488 79620
rect 131540 79568 131546 79620
rect 131822 79608 131850 79908
rect 132080 79840 132086 79892
rect 132138 79880 132144 79892
rect 132138 79840 132172 79880
rect 131988 79772 131994 79824
rect 132046 79772 132052 79824
rect 132006 79688 132034 79772
rect 132144 79688 132172 79840
rect 132282 79756 132310 79908
rect 132218 79704 132224 79756
rect 132276 79716 132310 79756
rect 132276 79704 132282 79716
rect 132374 79688 132402 79908
rect 132632 79880 132638 79892
rect 132604 79840 132638 79880
rect 132690 79840 132696 79892
rect 132724 79840 132730 79892
rect 132782 79840 132788 79892
rect 132604 79756 132632 79840
rect 132586 79704 132592 79756
rect 132644 79704 132650 79756
rect 132742 79688 132770 79840
rect 132006 79648 132040 79688
rect 132034 79636 132040 79648
rect 132092 79636 132098 79688
rect 132126 79636 132132 79688
rect 132184 79636 132190 79688
rect 132310 79636 132316 79688
rect 132368 79648 132402 79688
rect 132368 79636 132374 79648
rect 132678 79636 132684 79688
rect 132736 79648 132770 79688
rect 132736 79636 132742 79648
rect 133018 79620 133046 79920
rect 133184 79908 133190 79920
rect 133242 79908 133248 79960
rect 133644 79908 133650 79960
rect 133702 79908 133708 79960
rect 133092 79840 133098 79892
rect 133150 79880 133156 79892
rect 133150 79840 133184 79880
rect 133460 79840 133466 79892
rect 133518 79840 133524 79892
rect 133156 79756 133184 79840
rect 133138 79704 133144 79756
rect 133196 79704 133202 79756
rect 131942 79608 131948 79620
rect 131822 79580 131948 79608
rect 131942 79568 131948 79580
rect 132000 79568 132006 79620
rect 133018 79580 133052 79620
rect 133046 79568 133052 79580
rect 133104 79568 133110 79620
rect 132678 79500 132684 79552
rect 132736 79540 132742 79552
rect 133478 79540 133506 79840
rect 133662 79688 133690 79908
rect 133598 79636 133604 79688
rect 133656 79648 133690 79688
rect 133656 79636 133662 79648
rect 132736 79512 133506 79540
rect 132736 79500 132742 79512
rect 130344 79376 130838 79404
rect 130344 79364 130350 79376
rect 133506 79364 133512 79416
rect 133564 79404 133570 79416
rect 133754 79404 133782 79988
rect 136606 79988 137186 80016
rect 136606 79960 136634 79988
rect 134012 79908 134018 79960
rect 134070 79908 134076 79960
rect 134564 79908 134570 79960
rect 134622 79908 134628 79960
rect 134840 79948 134846 79960
rect 134674 79920 134846 79948
rect 134030 79824 134058 79908
rect 134196 79840 134202 79892
rect 134254 79880 134260 79892
rect 134254 79840 134288 79880
rect 134380 79840 134386 79892
rect 134438 79840 134444 79892
rect 133966 79772 133972 79824
rect 134024 79784 134058 79824
rect 134024 79772 134030 79784
rect 134104 79772 134110 79824
rect 134162 79772 134168 79824
rect 134122 79676 134150 79772
rect 134076 79648 134150 79676
rect 134076 79620 134104 79648
rect 134260 79620 134288 79840
rect 134058 79568 134064 79620
rect 134116 79568 134122 79620
rect 134242 79568 134248 79620
rect 134300 79568 134306 79620
rect 134150 79500 134156 79552
rect 134208 79540 134214 79552
rect 134398 79540 134426 79840
rect 134582 79812 134610 79908
rect 134536 79784 134610 79812
rect 134536 79756 134564 79784
rect 134518 79704 134524 79756
rect 134576 79704 134582 79756
rect 134674 79744 134702 79920
rect 134840 79908 134846 79920
rect 134898 79908 134904 79960
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 135484 79908 135490 79960
rect 135542 79908 135548 79960
rect 135576 79908 135582 79960
rect 135634 79908 135640 79960
rect 135852 79908 135858 79960
rect 135910 79908 135916 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 136312 79908 136318 79960
rect 136370 79908 136376 79960
rect 136404 79908 136410 79960
rect 136462 79908 136468 79960
rect 136588 79908 136594 79960
rect 136646 79908 136652 79960
rect 137048 79908 137054 79960
rect 137106 79908 137112 79960
rect 135024 79840 135030 79892
rect 135082 79840 135088 79892
rect 135042 79812 135070 79840
rect 134628 79716 134702 79744
rect 134858 79784 135070 79812
rect 134628 79688 134656 79716
rect 134610 79636 134616 79688
rect 134668 79636 134674 79688
rect 134702 79636 134708 79688
rect 134760 79676 134766 79688
rect 134858 79676 134886 79784
rect 135226 79744 135254 79908
rect 135300 79840 135306 79892
rect 135358 79880 135364 79892
rect 135358 79840 135392 79880
rect 135364 79756 135392 79840
rect 135502 79756 135530 79908
rect 134760 79648 134886 79676
rect 135088 79716 135254 79744
rect 134760 79636 134766 79648
rect 135088 79620 135116 79716
rect 135346 79704 135352 79756
rect 135404 79704 135410 79756
rect 135438 79704 135444 79756
rect 135496 79716 135530 79756
rect 135496 79704 135502 79716
rect 135070 79568 135076 79620
rect 135128 79568 135134 79620
rect 135254 79568 135260 79620
rect 135312 79608 135318 79620
rect 135594 79608 135622 79908
rect 135760 79772 135766 79824
rect 135818 79772 135824 79824
rect 135778 79688 135806 79772
rect 135714 79636 135720 79688
rect 135772 79648 135806 79688
rect 135870 79688 135898 79908
rect 136036 79840 136042 79892
rect 136094 79840 136100 79892
rect 136238 79880 136266 79908
rect 136192 79852 136266 79880
rect 135870 79648 135904 79688
rect 135772 79636 135778 79648
rect 135898 79636 135904 79648
rect 135956 79636 135962 79688
rect 135312 79580 135622 79608
rect 135312 79568 135318 79580
rect 134208 79512 134426 79540
rect 134208 79500 134214 79512
rect 135622 79500 135628 79552
rect 135680 79540 135686 79552
rect 136054 79540 136082 79840
rect 136192 79688 136220 79852
rect 136330 79812 136358 79908
rect 136284 79784 136358 79812
rect 136284 79688 136312 79784
rect 136422 79756 136450 79908
rect 137066 79880 137094 79908
rect 136790 79852 137094 79880
rect 136680 79772 136686 79824
rect 136738 79772 136744 79824
rect 136358 79704 136364 79756
rect 136416 79716 136450 79756
rect 136416 79704 136422 79716
rect 136174 79636 136180 79688
rect 136232 79636 136238 79688
rect 136266 79636 136272 79688
rect 136324 79636 136330 79688
rect 135680 79512 136082 79540
rect 135680 79500 135686 79512
rect 136698 79472 136726 79772
rect 136790 79688 136818 79852
rect 137158 79812 137186 79988
rect 137710 79960 137738 80056
rect 139320 79988 139946 80016
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137692 79908 137698 79960
rect 137750 79908 137756 79960
rect 137968 79908 137974 79960
rect 138026 79948 138032 79960
rect 138026 79920 138152 79948
rect 138026 79908 138032 79920
rect 137324 79840 137330 79892
rect 137382 79840 137388 79892
rect 137020 79784 137186 79812
rect 136790 79648 136824 79688
rect 136818 79636 136824 79648
rect 136876 79636 136882 79688
rect 136818 79500 136824 79552
rect 136876 79540 136882 79552
rect 137020 79540 137048 79784
rect 137342 79688 137370 79840
rect 137278 79636 137284 79688
rect 137336 79648 137370 79688
rect 137336 79636 137342 79648
rect 136876 79512 137048 79540
rect 137618 79552 137646 79908
rect 137784 79840 137790 79892
rect 137842 79880 137848 79892
rect 137842 79852 138060 79880
rect 137842 79840 137848 79852
rect 137618 79512 137652 79552
rect 136876 79500 136882 79512
rect 137646 79500 137652 79512
rect 137704 79500 137710 79552
rect 137738 79500 137744 79552
rect 137796 79540 137802 79552
rect 138032 79540 138060 79852
rect 138124 79620 138152 79920
rect 138244 79908 138250 79960
rect 138302 79908 138308 79960
rect 138336 79908 138342 79960
rect 138394 79908 138400 79960
rect 138520 79948 138526 79960
rect 138492 79908 138526 79948
rect 138578 79908 138584 79960
rect 138612 79908 138618 79960
rect 138670 79908 138676 79960
rect 138704 79908 138710 79960
rect 138762 79908 138768 79960
rect 138980 79908 138986 79960
rect 139038 79908 139044 79960
rect 139164 79948 139170 79960
rect 139136 79908 139170 79948
rect 139222 79908 139228 79960
rect 138262 79620 138290 79908
rect 138354 79688 138382 79908
rect 138492 79688 138520 79908
rect 138630 79880 138658 79908
rect 138584 79852 138658 79880
rect 138354 79648 138388 79688
rect 138382 79636 138388 79648
rect 138440 79636 138446 79688
rect 138474 79636 138480 79688
rect 138532 79636 138538 79688
rect 138106 79568 138112 79620
rect 138164 79568 138170 79620
rect 138262 79580 138296 79620
rect 138290 79568 138296 79580
rect 138348 79568 138354 79620
rect 137796 79512 138060 79540
rect 138584 79540 138612 79852
rect 138722 79812 138750 79908
rect 138796 79840 138802 79892
rect 138854 79840 138860 79892
rect 138888 79840 138894 79892
rect 138946 79840 138952 79892
rect 138676 79784 138750 79812
rect 138676 79756 138704 79784
rect 138814 79756 138842 79840
rect 138658 79704 138664 79756
rect 138716 79704 138722 79756
rect 138750 79704 138756 79756
rect 138808 79716 138842 79756
rect 138906 79756 138934 79840
rect 138998 79812 139026 79908
rect 139136 79824 139164 79908
rect 138998 79784 139072 79812
rect 139044 79756 139072 79784
rect 139118 79772 139124 79824
rect 139176 79772 139182 79824
rect 138906 79716 138940 79756
rect 138808 79704 138814 79716
rect 138934 79704 138940 79716
rect 138992 79704 138998 79756
rect 139026 79704 139032 79756
rect 139084 79704 139090 79756
rect 139026 79540 139032 79552
rect 138584 79512 139032 79540
rect 137796 79500 137802 79512
rect 139026 79500 139032 79512
rect 139084 79500 139090 79552
rect 139320 79540 139348 79988
rect 139918 79960 139946 79988
rect 139624 79908 139630 79960
rect 139682 79908 139688 79960
rect 139716 79908 139722 79960
rect 139774 79908 139780 79960
rect 139808 79908 139814 79960
rect 139866 79908 139872 79960
rect 139900 79908 139906 79960
rect 139958 79908 139964 79960
rect 139992 79908 139998 79960
rect 140050 79908 140056 79960
rect 140176 79908 140182 79960
rect 140234 79908 140240 79960
rect 140268 79908 140274 79960
rect 140326 79908 140332 79960
rect 140360 79908 140366 79960
rect 140418 79908 140424 79960
rect 140452 79908 140458 79960
rect 140510 79948 140516 79960
rect 141464 79948 141470 79960
rect 140510 79920 140958 79948
rect 140510 79908 140516 79920
rect 139532 79880 139538 79892
rect 139504 79840 139538 79880
rect 139590 79840 139596 79892
rect 139504 79676 139532 79840
rect 139642 79812 139670 79908
rect 139596 79784 139670 79812
rect 139596 79756 139624 79784
rect 139734 79756 139762 79908
rect 139826 79880 139854 79908
rect 139826 79852 139946 79880
rect 139918 79756 139946 79852
rect 139578 79704 139584 79756
rect 139636 79704 139642 79756
rect 139670 79704 139676 79756
rect 139728 79716 139762 79756
rect 139728 79704 139734 79716
rect 139854 79704 139860 79756
rect 139912 79716 139946 79756
rect 139912 79704 139918 79716
rect 139762 79676 139768 79688
rect 139504 79648 139768 79676
rect 139762 79636 139768 79648
rect 139820 79636 139826 79688
rect 140010 79676 140038 79908
rect 140194 79880 140222 79908
rect 140148 79852 140222 79880
rect 140148 79756 140176 79852
rect 140286 79824 140314 79908
rect 140222 79772 140228 79824
rect 140280 79784 140314 79824
rect 140378 79824 140406 79908
rect 140820 79840 140826 79892
rect 140878 79840 140884 79892
rect 140378 79784 140412 79824
rect 140280 79772 140286 79784
rect 140406 79772 140412 79784
rect 140464 79772 140470 79824
rect 140130 79704 140136 79756
rect 140188 79704 140194 79756
rect 140838 79744 140866 79840
rect 140792 79716 140866 79744
rect 140314 79676 140320 79688
rect 140010 79648 140320 79676
rect 140314 79636 140320 79648
rect 140372 79636 140378 79688
rect 139578 79540 139584 79552
rect 139320 79512 139584 79540
rect 139578 79500 139584 79512
rect 139636 79500 139642 79552
rect 140792 79540 140820 79716
rect 140930 79688 140958 79920
rect 141252 79920 141470 79948
rect 141096 79772 141102 79824
rect 141154 79812 141160 79824
rect 141154 79772 141188 79812
rect 141160 79688 141188 79772
rect 140866 79636 140872 79688
rect 140924 79648 140958 79688
rect 140924 79636 140930 79648
rect 141142 79636 141148 79688
rect 141200 79636 141206 79688
rect 141252 79620 141280 79920
rect 141464 79908 141470 79920
rect 141522 79908 141528 79960
rect 141648 79908 141654 79960
rect 141706 79908 141712 79960
rect 141740 79908 141746 79960
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141666 79880 141694 79908
rect 141528 79852 141694 79880
rect 141234 79568 141240 79620
rect 141292 79568 141298 79620
rect 141050 79540 141056 79552
rect 140792 79512 141056 79540
rect 141050 79500 141056 79512
rect 141108 79500 141114 79552
rect 138842 79472 138848 79484
rect 136698 79444 138848 79472
rect 138842 79432 138848 79444
rect 138900 79432 138906 79484
rect 140958 79432 140964 79484
rect 141016 79472 141022 79484
rect 141528 79472 141556 79852
rect 141758 79824 141786 79908
rect 141694 79772 141700 79824
rect 141752 79784 141786 79824
rect 141752 79772 141758 79784
rect 141850 79756 141878 79908
rect 142016 79880 142022 79892
rect 141988 79840 142022 79880
rect 142074 79840 142080 79892
rect 141850 79716 141884 79756
rect 141878 79704 141884 79716
rect 141936 79704 141942 79756
rect 141786 79636 141792 79688
rect 141844 79676 141850 79688
rect 141988 79676 142016 79840
rect 142126 79812 142154 80056
rect 144886 79988 145834 80016
rect 144886 79960 144914 79988
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 142292 79908 142298 79960
rect 142350 79908 142356 79960
rect 143488 79908 143494 79960
rect 143546 79908 143552 79960
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 144960 79908 144966 79960
rect 145018 79908 145024 79960
rect 145052 79908 145058 79960
rect 145110 79908 145116 79960
rect 145144 79908 145150 79960
rect 145202 79908 145208 79960
rect 145236 79908 145242 79960
rect 145294 79908 145300 79960
rect 145604 79948 145610 79960
rect 145530 79920 145610 79948
rect 142080 79784 142154 79812
rect 142080 79756 142108 79784
rect 142062 79704 142068 79756
rect 142120 79704 142126 79756
rect 141844 79648 142016 79676
rect 141844 79636 141850 79648
rect 141016 79444 141556 79472
rect 141016 79432 141022 79444
rect 142218 79404 142246 79908
rect 142310 79472 142338 79908
rect 142660 79840 142666 79892
rect 142718 79840 142724 79892
rect 142752 79840 142758 79892
rect 142810 79840 142816 79892
rect 143212 79840 143218 79892
rect 143270 79840 143276 79892
rect 142678 79620 142706 79840
rect 142770 79744 142798 79840
rect 142770 79716 142936 79744
rect 142908 79620 142936 79716
rect 143230 79688 143258 79840
rect 143506 79824 143534 79908
rect 143580 79840 143586 79892
rect 143638 79840 143644 79892
rect 143764 79840 143770 79892
rect 143822 79840 143828 79892
rect 144040 79840 144046 79892
rect 144098 79880 144104 79892
rect 144098 79840 144132 79880
rect 144316 79840 144322 79892
rect 144374 79880 144380 79892
rect 144978 79880 145006 79908
rect 144374 79852 144730 79880
rect 144374 79840 144380 79852
rect 143442 79772 143448 79824
rect 143500 79784 143534 79824
rect 143500 79772 143506 79784
rect 143598 79688 143626 79840
rect 143672 79772 143678 79824
rect 143730 79772 143736 79824
rect 143230 79648 143264 79688
rect 143258 79636 143264 79648
rect 143316 79636 143322 79688
rect 143534 79636 143540 79688
rect 143592 79648 143626 79688
rect 143592 79636 143598 79648
rect 142678 79580 142712 79620
rect 142706 79568 142712 79580
rect 142764 79568 142770 79620
rect 142890 79568 142896 79620
rect 142948 79568 142954 79620
rect 143690 79540 143718 79772
rect 143782 79608 143810 79840
rect 143948 79772 143954 79824
rect 144006 79772 144012 79824
rect 143966 79688 143994 79772
rect 144104 79756 144132 79840
rect 144086 79704 144092 79756
rect 144144 79704 144150 79756
rect 143902 79636 143908 79688
rect 143960 79648 143994 79688
rect 143960 79636 143966 79648
rect 144702 79620 144730 79852
rect 144932 79852 145006 79880
rect 144776 79772 144782 79824
rect 144834 79772 144840 79824
rect 144794 79744 144822 79772
rect 144932 79756 144960 79852
rect 145070 79756 145098 79908
rect 144794 79716 144868 79744
rect 144840 79620 144868 79716
rect 144914 79704 144920 79756
rect 144972 79704 144978 79756
rect 145006 79704 145012 79756
rect 145064 79716 145098 79756
rect 145064 79704 145070 79716
rect 144270 79608 144276 79620
rect 143782 79580 144276 79608
rect 144270 79568 144276 79580
rect 144328 79568 144334 79620
rect 144702 79580 144736 79620
rect 144730 79568 144736 79580
rect 144788 79568 144794 79620
rect 144822 79568 144828 79620
rect 144880 79568 144886 79620
rect 145162 79608 145190 79908
rect 144932 79580 145190 79608
rect 143994 79540 144000 79552
rect 143690 79512 144000 79540
rect 143994 79500 144000 79512
rect 144052 79500 144058 79552
rect 144546 79500 144552 79552
rect 144604 79540 144610 79552
rect 144932 79540 144960 79580
rect 144604 79512 144960 79540
rect 144604 79500 144610 79512
rect 145006 79500 145012 79552
rect 145064 79540 145070 79552
rect 145254 79540 145282 79908
rect 145420 79772 145426 79824
rect 145478 79772 145484 79824
rect 145438 79744 145466 79772
rect 145392 79716 145466 79744
rect 145392 79620 145420 79716
rect 145530 79620 145558 79920
rect 145604 79908 145610 79920
rect 145662 79908 145668 79960
rect 145696 79908 145702 79960
rect 145754 79908 145760 79960
rect 145714 79824 145742 79908
rect 145650 79772 145656 79824
rect 145708 79784 145742 79824
rect 145708 79772 145714 79784
rect 145806 79620 145834 79988
rect 145898 79960 145926 80124
rect 145880 79908 145886 79960
rect 145938 79908 145944 79960
rect 146156 79908 146162 79960
rect 146214 79908 146220 79960
rect 146432 79908 146438 79960
rect 146490 79908 146496 79960
rect 146616 79908 146622 79960
rect 146674 79908 146680 79960
rect 146708 79908 146714 79960
rect 146766 79908 146772 79960
rect 147168 79908 147174 79960
rect 147226 79908 147232 79960
rect 147260 79908 147266 79960
rect 147318 79908 147324 79960
rect 147444 79908 147450 79960
rect 147502 79908 147508 79960
rect 147904 79908 147910 79960
rect 147962 79908 147968 79960
rect 148272 79908 148278 79960
rect 148330 79908 148336 79960
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 149836 79948 149842 79960
rect 149808 79908 149842 79948
rect 149894 79908 149900 79960
rect 149928 79908 149934 79960
rect 149986 79908 149992 79960
rect 150020 79908 150026 79960
rect 150078 79908 150084 79960
rect 150112 79908 150118 79960
rect 150170 79908 150176 79960
rect 145972 79840 145978 79892
rect 146030 79840 146036 79892
rect 145990 79756 146018 79840
rect 145926 79704 145932 79756
rect 145984 79716 146018 79756
rect 145984 79704 145990 79716
rect 146018 79636 146024 79688
rect 146076 79676 146082 79688
rect 146174 79676 146202 79908
rect 146076 79648 146202 79676
rect 146076 79636 146082 79648
rect 145374 79568 145380 79620
rect 145432 79568 145438 79620
rect 145466 79568 145472 79620
rect 145524 79580 145558 79620
rect 145524 79568 145530 79580
rect 145742 79568 145748 79620
rect 145800 79580 145834 79620
rect 146450 79620 146478 79908
rect 146450 79580 146484 79620
rect 145800 79568 145806 79580
rect 146478 79568 146484 79580
rect 146536 79568 146542 79620
rect 145064 79512 145282 79540
rect 145064 79500 145070 79512
rect 146386 79500 146392 79552
rect 146444 79540 146450 79552
rect 146634 79540 146662 79908
rect 146726 79620 146754 79908
rect 146892 79840 146898 79892
rect 146950 79840 146956 79892
rect 147076 79880 147082 79892
rect 147002 79852 147082 79880
rect 146910 79688 146938 79840
rect 146846 79636 146852 79688
rect 146904 79648 146938 79688
rect 146904 79636 146910 79648
rect 147002 79620 147030 79852
rect 147076 79840 147082 79852
rect 147134 79840 147140 79892
rect 147186 79812 147214 79908
rect 147094 79784 147214 79812
rect 147278 79824 147306 79908
rect 147278 79784 147312 79824
rect 147094 79676 147122 79784
rect 147306 79772 147312 79784
rect 147364 79772 147370 79824
rect 147462 79812 147490 79908
rect 147628 79840 147634 79892
rect 147686 79840 147692 79892
rect 147462 79784 147536 79812
rect 147508 79688 147536 79784
rect 147214 79676 147220 79688
rect 147094 79648 147220 79676
rect 147214 79636 147220 79648
rect 147272 79636 147278 79688
rect 147490 79636 147496 79688
rect 147548 79636 147554 79688
rect 146726 79580 146760 79620
rect 146754 79568 146760 79580
rect 146812 79568 146818 79620
rect 146938 79568 146944 79620
rect 146996 79580 147030 79620
rect 146996 79568 147002 79580
rect 146444 79512 146662 79540
rect 146444 79500 146450 79512
rect 142614 79472 142620 79484
rect 142310 79444 142620 79472
rect 142614 79432 142620 79444
rect 142672 79432 142678 79484
rect 143810 79432 143816 79484
rect 143868 79472 143874 79484
rect 147646 79472 147674 79840
rect 143868 79444 147674 79472
rect 147922 79484 147950 79908
rect 148290 79824 148318 79908
rect 148916 79840 148922 79892
rect 148974 79840 148980 79892
rect 148180 79772 148186 79824
rect 148238 79772 148244 79824
rect 148290 79784 148324 79824
rect 148318 79772 148324 79784
rect 148376 79772 148382 79824
rect 148198 79688 148226 79772
rect 148198 79648 148232 79688
rect 148226 79636 148232 79648
rect 148284 79636 148290 79688
rect 148686 79500 148692 79552
rect 148744 79540 148750 79552
rect 148934 79540 148962 79840
rect 149210 79744 149238 79908
rect 149652 79880 149658 79892
rect 149532 79852 149658 79880
rect 149284 79772 149290 79824
rect 149342 79772 149348 79824
rect 149164 79716 149238 79744
rect 149164 79552 149192 79716
rect 149302 79620 149330 79772
rect 149238 79568 149244 79620
rect 149296 79580 149330 79620
rect 149296 79568 149302 79580
rect 148744 79512 148962 79540
rect 148744 79500 148750 79512
rect 149146 79500 149152 79552
rect 149204 79500 149210 79552
rect 149330 79500 149336 79552
rect 149388 79540 149394 79552
rect 149532 79540 149560 79852
rect 149652 79840 149658 79852
rect 149710 79840 149716 79892
rect 149808 79688 149836 79908
rect 149946 79880 149974 79908
rect 149900 79852 149974 79880
rect 149900 79756 149928 79852
rect 150038 79812 150066 79908
rect 149992 79784 150066 79812
rect 149992 79756 150020 79784
rect 150130 79756 150158 79908
rect 149882 79704 149888 79756
rect 149940 79704 149946 79756
rect 149974 79704 149980 79756
rect 150032 79704 150038 79756
rect 150066 79704 150072 79756
rect 150124 79716 150158 79756
rect 150124 79704 150130 79716
rect 149790 79636 149796 79688
rect 149848 79636 149854 79688
rect 150158 79568 150164 79620
rect 150216 79608 150222 79620
rect 150360 79608 150388 80124
rect 150958 79988 151170 80016
rect 150958 79960 150986 79988
rect 150480 79908 150486 79960
rect 150538 79908 150544 79960
rect 150572 79908 150578 79960
rect 150630 79908 150636 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 150940 79908 150946 79960
rect 150998 79908 151004 79960
rect 150216 79580 150388 79608
rect 150216 79568 150222 79580
rect 150498 79552 150526 79908
rect 150590 79744 150618 79908
rect 150774 79824 150802 79908
rect 151032 79840 151038 79892
rect 151090 79840 151096 79892
rect 150774 79784 150808 79824
rect 150802 79772 150808 79784
rect 150860 79772 150866 79824
rect 150894 79744 150900 79756
rect 150590 79716 150900 79744
rect 150894 79704 150900 79716
rect 150952 79704 150958 79756
rect 150710 79636 150716 79688
rect 150768 79676 150774 79688
rect 151050 79676 151078 79840
rect 150768 79648 151078 79676
rect 150768 79636 150774 79648
rect 150986 79568 150992 79620
rect 151044 79608 151050 79620
rect 151142 79608 151170 79988
rect 151832 79988 152458 80016
rect 151400 79908 151406 79960
rect 151458 79908 151464 79960
rect 151308 79840 151314 79892
rect 151366 79840 151372 79892
rect 151044 79580 151170 79608
rect 151044 79568 151050 79580
rect 151326 79552 151354 79840
rect 151418 79756 151446 79908
rect 151418 79716 151452 79756
rect 151446 79704 151452 79716
rect 151504 79704 151510 79756
rect 151832 79552 151860 79988
rect 152430 79960 152458 79988
rect 152136 79908 152142 79960
rect 152194 79948 152200 79960
rect 152194 79920 152366 79948
rect 152194 79908 152200 79920
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 151998 79568 152004 79620
rect 152056 79608 152062 79620
rect 152246 79608 152274 79840
rect 152056 79580 152274 79608
rect 152056 79568 152062 79580
rect 152338 79552 152366 79920
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 153166 79880 153194 80192
rect 154546 80016 154574 80328
rect 177022 80316 177028 80368
rect 177080 80356 177086 80368
rect 186286 80356 186314 80668
rect 580534 80656 580540 80668
rect 580592 80656 580598 80708
rect 177080 80328 186314 80356
rect 177080 80316 177086 80328
rect 153258 79988 154574 80016
rect 154638 80260 171686 80288
rect 153258 79960 153286 79988
rect 154638 79960 154666 80260
rect 158686 80192 163728 80220
rect 158686 80084 158714 80192
rect 163700 80152 163728 80192
rect 163884 80192 170766 80220
rect 163884 80152 163912 80192
rect 163700 80124 163912 80152
rect 164206 80124 165062 80152
rect 164206 80084 164234 80124
rect 158686 80056 158806 80084
rect 158778 79960 158806 80056
rect 160664 80056 162026 80084
rect 160664 80016 160692 80056
rect 159146 79988 160692 80016
rect 159146 79960 159174 79988
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153700 79948 153706 79960
rect 153672 79908 153706 79948
rect 153758 79908 153764 79960
rect 153884 79908 153890 79960
rect 153942 79908 153948 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 155816 79908 155822 79960
rect 155874 79908 155880 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156000 79908 156006 79960
rect 156058 79908 156064 79960
rect 156092 79908 156098 79960
rect 156150 79908 156156 79960
rect 156460 79908 156466 79960
rect 156518 79908 156524 79960
rect 156736 79908 156742 79960
rect 156794 79948 156800 79960
rect 156794 79908 156828 79948
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 157012 79908 157018 79960
rect 157070 79908 157076 79960
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157748 79948 157754 79960
rect 157352 79920 157754 79948
rect 153166 79852 153240 79880
rect 153212 79824 153240 79852
rect 153424 79840 153430 79892
rect 153482 79840 153488 79892
rect 152780 79772 152786 79824
rect 152838 79772 152844 79824
rect 153194 79772 153200 79824
rect 153252 79772 153258 79824
rect 152798 79688 152826 79772
rect 153442 79688 153470 79840
rect 152734 79636 152740 79688
rect 152792 79648 152826 79688
rect 152792 79636 152798 79648
rect 153378 79636 153384 79688
rect 153436 79648 153470 79688
rect 153436 79636 153442 79648
rect 149388 79512 149560 79540
rect 149388 79500 149394 79512
rect 150434 79500 150440 79552
rect 150492 79512 150526 79552
rect 150492 79500 150498 79512
rect 151262 79500 151268 79552
rect 151320 79512 151354 79552
rect 151320 79500 151326 79512
rect 151814 79500 151820 79552
rect 151872 79500 151878 79552
rect 152274 79500 152280 79552
rect 152332 79512 152366 79552
rect 153672 79540 153700 79908
rect 153792 79880 153798 79892
rect 153764 79840 153798 79880
rect 153850 79840 153856 79892
rect 153764 79756 153792 79840
rect 153902 79756 153930 79908
rect 154160 79840 154166 79892
rect 154218 79840 154224 79892
rect 153746 79704 153752 79756
rect 153804 79704 153810 79756
rect 153838 79704 153844 79756
rect 153896 79716 153930 79756
rect 154178 79756 154206 79840
rect 154270 79812 154298 79908
rect 154896 79840 154902 79892
rect 154954 79840 154960 79892
rect 155172 79840 155178 79892
rect 155230 79840 155236 79892
rect 155448 79840 155454 79892
rect 155506 79840 155512 79892
rect 155834 79880 155862 79908
rect 155788 79852 155862 79880
rect 154270 79784 154528 79812
rect 154178 79716 154212 79756
rect 153896 79704 153902 79716
rect 154206 79704 154212 79716
rect 154264 79704 154270 79756
rect 154500 79688 154528 79784
rect 154482 79636 154488 79688
rect 154540 79636 154546 79688
rect 154574 79636 154580 79688
rect 154632 79676 154638 79688
rect 154914 79676 154942 79840
rect 154632 79648 154942 79676
rect 154632 79636 154638 79648
rect 154758 79568 154764 79620
rect 154816 79608 154822 79620
rect 155190 79608 155218 79840
rect 155466 79812 155494 79840
rect 155328 79784 155494 79812
rect 155328 79620 155356 79784
rect 155788 79756 155816 79852
rect 155926 79812 155954 79908
rect 155880 79784 155954 79812
rect 155880 79756 155908 79784
rect 155402 79704 155408 79756
rect 155460 79704 155466 79756
rect 155770 79704 155776 79756
rect 155828 79704 155834 79756
rect 155862 79704 155868 79756
rect 155920 79704 155926 79756
rect 156018 79744 156046 79908
rect 155972 79716 156046 79744
rect 154816 79580 155218 79608
rect 154816 79568 154822 79580
rect 155310 79568 155316 79620
rect 155368 79568 155374 79620
rect 154022 79540 154028 79552
rect 153672 79512 154028 79540
rect 152332 79500 152338 79512
rect 154022 79500 154028 79512
rect 154080 79500 154086 79552
rect 155420 79540 155448 79704
rect 155494 79540 155500 79552
rect 155420 79512 155500 79540
rect 155494 79500 155500 79512
rect 155552 79500 155558 79552
rect 155972 79540 156000 79716
rect 156110 79620 156138 79908
rect 156276 79840 156282 79892
rect 156334 79880 156340 79892
rect 156334 79840 156368 79880
rect 156340 79688 156368 79840
rect 156478 79744 156506 79908
rect 156552 79840 156558 79892
rect 156610 79840 156616 79892
rect 156644 79840 156650 79892
rect 156702 79840 156708 79892
rect 156432 79716 156506 79744
rect 156432 79688 156460 79716
rect 156570 79688 156598 79840
rect 156322 79636 156328 79688
rect 156380 79636 156386 79688
rect 156414 79636 156420 79688
rect 156472 79636 156478 79688
rect 156506 79636 156512 79688
rect 156564 79648 156598 79688
rect 156662 79688 156690 79840
rect 156800 79688 156828 79908
rect 156662 79648 156696 79688
rect 156564 79636 156570 79648
rect 156690 79636 156696 79648
rect 156748 79636 156754 79688
rect 156782 79636 156788 79688
rect 156840 79636 156846 79688
rect 156046 79568 156052 79620
rect 156104 79580 156138 79620
rect 156104 79568 156110 79580
rect 156230 79540 156236 79552
rect 155972 79512 156236 79540
rect 156230 79500 156236 79512
rect 156288 79500 156294 79552
rect 156938 79540 156966 79908
rect 157030 79620 157058 79908
rect 157214 79824 157242 79908
rect 157150 79772 157156 79824
rect 157208 79784 157242 79824
rect 157208 79772 157214 79784
rect 157030 79580 157064 79620
rect 157058 79568 157064 79580
rect 157116 79568 157122 79620
rect 157150 79540 157156 79552
rect 156938 79512 157156 79540
rect 157150 79500 157156 79512
rect 157208 79500 157214 79552
rect 157242 79500 157248 79552
rect 157300 79540 157306 79552
rect 157352 79540 157380 79920
rect 157748 79908 157754 79920
rect 157806 79908 157812 79960
rect 158392 79908 158398 79960
rect 158450 79908 158456 79960
rect 158668 79908 158674 79960
rect 158726 79908 158732 79960
rect 158760 79908 158766 79960
rect 158818 79908 158824 79960
rect 159128 79908 159134 79960
rect 159186 79908 159192 79960
rect 159864 79908 159870 79960
rect 159922 79908 159928 79960
rect 159956 79908 159962 79960
rect 160014 79908 160020 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160508 79908 160514 79960
rect 160566 79908 160572 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160968 79908 160974 79960
rect 161026 79908 161032 79960
rect 161244 79948 161250 79960
rect 161078 79920 161250 79948
rect 157472 79840 157478 79892
rect 157530 79840 157536 79892
rect 157656 79840 157662 79892
rect 157714 79840 157720 79892
rect 157840 79840 157846 79892
rect 157898 79840 157904 79892
rect 157300 79512 157380 79540
rect 157490 79552 157518 79840
rect 157674 79620 157702 79840
rect 157610 79568 157616 79620
rect 157668 79580 157702 79620
rect 157858 79620 157886 79840
rect 158208 79772 158214 79824
rect 158266 79772 158272 79824
rect 158226 79688 158254 79772
rect 158410 79756 158438 79908
rect 158484 79840 158490 79892
rect 158542 79880 158548 79892
rect 158542 79840 158576 79880
rect 158410 79716 158444 79756
rect 158438 79704 158444 79716
rect 158496 79704 158502 79756
rect 158162 79636 158168 79688
rect 158220 79648 158254 79688
rect 158220 79636 158226 79648
rect 157858 79580 157892 79620
rect 157668 79568 157674 79580
rect 157886 79568 157892 79580
rect 157944 79568 157950 79620
rect 158346 79568 158352 79620
rect 158404 79608 158410 79620
rect 158548 79608 158576 79840
rect 158686 79744 158714 79908
rect 158852 79840 158858 79892
rect 158910 79880 158916 79892
rect 158910 79852 158990 79880
rect 158910 79840 158916 79852
rect 158806 79744 158812 79756
rect 158686 79716 158812 79744
rect 158806 79704 158812 79716
rect 158864 79704 158870 79756
rect 158962 79676 158990 79852
rect 159036 79840 159042 79892
rect 159094 79840 159100 79892
rect 159220 79840 159226 79892
rect 159278 79840 159284 79892
rect 159404 79840 159410 79892
rect 159462 79880 159468 79892
rect 159588 79880 159594 79892
rect 159462 79840 159496 79880
rect 159054 79744 159082 79840
rect 159238 79812 159266 79840
rect 159238 79784 159404 79812
rect 159376 79756 159404 79784
rect 159054 79716 159220 79744
rect 159192 79688 159220 79716
rect 159358 79704 159364 79756
rect 159416 79704 159422 79756
rect 159082 79676 159088 79688
rect 158962 79648 159088 79676
rect 159082 79636 159088 79648
rect 159140 79636 159146 79688
rect 159174 79636 159180 79688
rect 159232 79636 159238 79688
rect 158404 79580 158576 79608
rect 158404 79568 158410 79580
rect 158990 79568 158996 79620
rect 159048 79608 159054 79620
rect 159468 79608 159496 79840
rect 159560 79840 159594 79880
rect 159646 79840 159652 79892
rect 159560 79756 159588 79840
rect 159542 79704 159548 79756
rect 159600 79704 159606 79756
rect 159048 79580 159496 79608
rect 159048 79568 159054 79580
rect 159882 79552 159910 79908
rect 159974 79676 160002 79908
rect 160048 79840 160054 79892
rect 160106 79840 160112 79892
rect 160066 79744 160094 79840
rect 160158 79812 160186 79908
rect 160158 79784 160324 79812
rect 160066 79716 160186 79744
rect 159974 79648 160048 79676
rect 160020 79620 160048 79648
rect 160158 79620 160186 79716
rect 160002 79568 160008 79620
rect 160060 79568 160066 79620
rect 160158 79580 160192 79620
rect 160186 79568 160192 79580
rect 160244 79568 160250 79620
rect 157490 79512 157524 79552
rect 157300 79500 157306 79512
rect 157518 79500 157524 79512
rect 157576 79500 157582 79552
rect 157702 79500 157708 79552
rect 157760 79540 157766 79552
rect 159634 79540 159640 79552
rect 157760 79512 159640 79540
rect 157760 79500 157766 79512
rect 159634 79500 159640 79512
rect 159692 79500 159698 79552
rect 159818 79500 159824 79552
rect 159876 79512 159910 79552
rect 159876 79500 159882 79512
rect 160094 79500 160100 79552
rect 160152 79540 160158 79552
rect 160296 79540 160324 79784
rect 160152 79512 160324 79540
rect 160152 79500 160158 79512
rect 160370 79500 160376 79552
rect 160428 79540 160434 79552
rect 160526 79540 160554 79908
rect 160618 79880 160646 79908
rect 160618 79852 160876 79880
rect 160692 79772 160698 79824
rect 160750 79812 160756 79824
rect 160750 79772 160784 79812
rect 160756 79608 160784 79772
rect 160848 79676 160876 79852
rect 160986 79824 161014 79908
rect 160922 79772 160928 79824
rect 160980 79784 161014 79824
rect 160980 79772 160986 79784
rect 161078 79688 161106 79920
rect 161244 79908 161250 79920
rect 161302 79908 161308 79960
rect 161520 79908 161526 79960
rect 161578 79908 161584 79960
rect 161796 79908 161802 79960
rect 161854 79908 161860 79960
rect 161152 79840 161158 79892
rect 161210 79840 161216 79892
rect 161170 79744 161198 79840
rect 161336 79772 161342 79824
rect 161394 79772 161400 79824
rect 161170 79716 161290 79744
rect 160922 79676 160928 79688
rect 160848 79648 160928 79676
rect 160922 79636 160928 79648
rect 160980 79636 160986 79688
rect 161078 79648 161112 79688
rect 161106 79636 161112 79648
rect 161164 79636 161170 79688
rect 161262 79620 161290 79716
rect 161354 79688 161382 79772
rect 161538 79756 161566 79908
rect 161814 79812 161842 79908
rect 161814 79784 161888 79812
rect 161538 79716 161572 79756
rect 161566 79704 161572 79716
rect 161624 79704 161630 79756
rect 161354 79648 161388 79688
rect 161382 79636 161388 79648
rect 161440 79636 161446 79688
rect 161014 79608 161020 79620
rect 160756 79580 161020 79608
rect 161014 79568 161020 79580
rect 161072 79568 161078 79620
rect 161262 79580 161296 79620
rect 161290 79568 161296 79580
rect 161348 79568 161354 79620
rect 160428 79512 160554 79540
rect 160428 79500 160434 79512
rect 147922 79444 147956 79484
rect 143868 79432 143874 79444
rect 147950 79432 147956 79444
rect 148008 79432 148014 79484
rect 148318 79432 148324 79484
rect 148376 79472 148382 79484
rect 148376 79444 161244 79472
rect 148376 79432 148382 79444
rect 143074 79404 143080 79416
rect 133564 79376 133782 79404
rect 133846 79376 136312 79404
rect 142218 79376 143080 79404
rect 133564 79364 133570 79376
rect 127894 79336 127900 79348
rect 123496 79308 127900 79336
rect 127894 79296 127900 79308
rect 127952 79296 127958 79348
rect 128722 79296 128728 79348
rect 128780 79336 128786 79348
rect 133846 79336 133874 79376
rect 128780 79308 133874 79336
rect 136284 79336 136312 79376
rect 143074 79364 143080 79376
rect 143132 79364 143138 79416
rect 143534 79364 143540 79416
rect 143592 79404 143598 79416
rect 161216 79404 161244 79444
rect 161750 79432 161756 79484
rect 161808 79472 161814 79484
rect 161860 79472 161888 79784
rect 161998 79540 162026 80056
rect 163102 80056 164234 80084
rect 162274 79988 162992 80016
rect 162274 79960 162302 79988
rect 162256 79908 162262 79960
rect 162314 79908 162320 79960
rect 162440 79908 162446 79960
rect 162498 79908 162504 79960
rect 162532 79908 162538 79960
rect 162590 79908 162596 79960
rect 162808 79908 162814 79960
rect 162866 79908 162872 79960
rect 162458 79824 162486 79908
rect 162072 79772 162078 79824
rect 162130 79772 162136 79824
rect 162164 79772 162170 79824
rect 162222 79772 162228 79824
rect 162348 79772 162354 79824
rect 162406 79772 162412 79824
rect 162440 79772 162446 79824
rect 162498 79772 162504 79824
rect 162090 79688 162118 79772
rect 162182 79744 162210 79772
rect 162182 79716 162256 79744
rect 162228 79688 162256 79716
rect 162366 79688 162394 79772
rect 162090 79648 162124 79688
rect 162118 79636 162124 79648
rect 162176 79636 162182 79688
rect 162210 79636 162216 79688
rect 162268 79636 162274 79688
rect 162302 79636 162308 79688
rect 162360 79648 162394 79688
rect 162360 79636 162366 79648
rect 162550 79620 162578 79908
rect 162624 79772 162630 79824
rect 162682 79772 162688 79824
rect 162642 79688 162670 79772
rect 162642 79648 162676 79688
rect 162670 79636 162676 79648
rect 162728 79636 162734 79688
rect 162486 79568 162492 79620
rect 162544 79580 162578 79620
rect 162544 79568 162550 79580
rect 162578 79540 162584 79552
rect 161998 79512 162584 79540
rect 162578 79500 162584 79512
rect 162636 79500 162642 79552
rect 162826 79540 162854 79908
rect 162964 79688 162992 79988
rect 163102 79960 163130 80056
rect 164160 79988 164970 80016
rect 163084 79908 163090 79960
rect 163142 79908 163148 79960
rect 163452 79908 163458 79960
rect 163510 79908 163516 79960
rect 163636 79908 163642 79960
rect 163694 79908 163700 79960
rect 163912 79908 163918 79960
rect 163970 79908 163976 79960
rect 164004 79908 164010 79960
rect 164062 79948 164068 79960
rect 164062 79908 164096 79948
rect 162946 79636 162952 79688
rect 163004 79636 163010 79688
rect 163470 79552 163498 79908
rect 162946 79540 162952 79552
rect 162826 79512 162952 79540
rect 162946 79500 162952 79512
rect 163004 79500 163010 79552
rect 163470 79512 163504 79552
rect 163498 79500 163504 79512
rect 163556 79500 163562 79552
rect 161808 79444 161888 79472
rect 161808 79432 161814 79444
rect 162670 79432 162676 79484
rect 162728 79472 162734 79484
rect 163130 79472 163136 79484
rect 162728 79444 163136 79472
rect 162728 79432 162734 79444
rect 163130 79432 163136 79444
rect 163188 79432 163194 79484
rect 163654 79472 163682 79908
rect 163820 79772 163826 79824
rect 163878 79772 163884 79824
rect 163838 79620 163866 79772
rect 163930 79688 163958 79908
rect 164068 79688 164096 79908
rect 163930 79648 163964 79688
rect 163958 79636 163964 79648
rect 164016 79636 164022 79688
rect 164050 79636 164056 79688
rect 164108 79636 164114 79688
rect 163838 79580 163872 79620
rect 163866 79568 163872 79580
rect 163924 79568 163930 79620
rect 163774 79472 163780 79484
rect 163654 79444 163780 79472
rect 163774 79432 163780 79444
rect 163832 79432 163838 79484
rect 164160 79472 164188 79988
rect 164942 79960 164970 79988
rect 164280 79948 164286 79960
rect 164252 79908 164286 79948
rect 164338 79908 164344 79960
rect 164648 79908 164654 79960
rect 164706 79908 164712 79960
rect 164832 79908 164838 79960
rect 164890 79908 164896 79960
rect 164924 79908 164930 79960
rect 164982 79908 164988 79960
rect 164252 79688 164280 79908
rect 164464 79840 164470 79892
rect 164522 79840 164528 79892
rect 164234 79636 164240 79688
rect 164292 79636 164298 79688
rect 164482 79540 164510 79840
rect 164666 79620 164694 79908
rect 164602 79568 164608 79620
rect 164660 79580 164694 79620
rect 164660 79568 164666 79580
rect 164694 79540 164700 79552
rect 164482 79512 164700 79540
rect 164694 79500 164700 79512
rect 164752 79500 164758 79552
rect 164510 79472 164516 79484
rect 164160 79444 164516 79472
rect 164510 79432 164516 79444
rect 164568 79432 164574 79484
rect 164850 79472 164878 79908
rect 165034 79824 165062 80124
rect 165954 79988 166442 80016
rect 165954 79960 165982 79988
rect 165568 79908 165574 79960
rect 165626 79908 165632 79960
rect 165660 79908 165666 79960
rect 165718 79908 165724 79960
rect 165936 79908 165942 79960
rect 165994 79908 166000 79960
rect 166304 79908 166310 79960
rect 166362 79908 166368 79960
rect 165292 79840 165298 79892
rect 165350 79840 165356 79892
rect 164970 79772 164976 79824
rect 165028 79784 165062 79824
rect 165028 79772 165034 79784
rect 165200 79772 165206 79824
rect 165258 79772 165264 79824
rect 165062 79744 165068 79756
rect 164988 79716 165068 79744
rect 164988 79688 165016 79716
rect 165062 79704 165068 79716
rect 165120 79704 165126 79756
rect 164970 79636 164976 79688
rect 165028 79636 165034 79688
rect 165218 79552 165246 79772
rect 165310 79620 165338 79840
rect 165586 79620 165614 79908
rect 165678 79676 165706 79908
rect 165752 79772 165758 79824
rect 165810 79812 165816 79824
rect 165982 79812 165988 79824
rect 165810 79784 165988 79812
rect 165810 79772 165816 79784
rect 165982 79772 165988 79784
rect 166040 79772 166046 79824
rect 165890 79704 165896 79756
rect 165948 79744 165954 79756
rect 165948 79716 166028 79744
rect 165948 79704 165954 79716
rect 165678 79648 165936 79676
rect 165908 79620 165936 79648
rect 165310 79580 165344 79620
rect 165338 79568 165344 79580
rect 165396 79568 165402 79620
rect 165586 79580 165620 79620
rect 165614 79568 165620 79580
rect 165672 79568 165678 79620
rect 165890 79568 165896 79620
rect 165948 79568 165954 79620
rect 165218 79512 165252 79552
rect 165246 79500 165252 79512
rect 165304 79500 165310 79552
rect 165798 79500 165804 79552
rect 165856 79540 165862 79552
rect 166000 79540 166028 79716
rect 165856 79512 166028 79540
rect 165856 79500 165862 79512
rect 165154 79472 165160 79484
rect 164850 79444 165160 79472
rect 165154 79432 165160 79444
rect 165212 79432 165218 79484
rect 165430 79432 165436 79484
rect 165488 79472 165494 79484
rect 166322 79472 166350 79908
rect 166414 79608 166442 79988
rect 166506 79988 166810 80016
rect 166506 79676 166534 79988
rect 166782 79960 166810 79988
rect 167610 79988 168098 80016
rect 167610 79960 167638 79988
rect 166580 79908 166586 79960
rect 166638 79908 166644 79960
rect 166672 79908 166678 79960
rect 166730 79908 166736 79960
rect 166764 79908 166770 79960
rect 166822 79908 166828 79960
rect 166856 79908 166862 79960
rect 166914 79908 166920 79960
rect 167408 79948 167414 79960
rect 167150 79920 167414 79948
rect 166598 79756 166626 79908
rect 166690 79812 166718 79908
rect 166690 79784 166764 79812
rect 166598 79716 166632 79756
rect 166626 79704 166632 79716
rect 166684 79704 166690 79756
rect 166506 79648 166672 79676
rect 166534 79608 166540 79620
rect 166414 79580 166540 79608
rect 166534 79568 166540 79580
rect 166592 79568 166598 79620
rect 165488 79444 166350 79472
rect 166644 79472 166672 79648
rect 166736 79540 166764 79784
rect 166874 79756 166902 79908
rect 166874 79716 166908 79756
rect 166902 79704 166908 79716
rect 166960 79704 166966 79756
rect 167150 79608 167178 79920
rect 167408 79908 167414 79920
rect 167466 79908 167472 79960
rect 167500 79908 167506 79960
rect 167558 79908 167564 79960
rect 167592 79908 167598 79960
rect 167650 79908 167656 79960
rect 167684 79908 167690 79960
rect 167742 79908 167748 79960
rect 167776 79908 167782 79960
rect 167834 79908 167840 79960
rect 167960 79908 167966 79960
rect 168018 79908 168024 79960
rect 167224 79840 167230 79892
rect 167282 79840 167288 79892
rect 167242 79676 167270 79840
rect 167518 79812 167546 79908
rect 167702 79812 167730 79908
rect 167518 79784 167592 79812
rect 167454 79676 167460 79688
rect 167242 79648 167460 79676
rect 167454 79636 167460 79648
rect 167512 79636 167518 79688
rect 167270 79608 167276 79620
rect 167150 79580 167276 79608
rect 167270 79568 167276 79580
rect 167328 79568 167334 79620
rect 167362 79568 167368 79620
rect 167420 79608 167426 79620
rect 167564 79608 167592 79784
rect 167656 79784 167730 79812
rect 167656 79756 167684 79784
rect 167794 79756 167822 79908
rect 167868 79840 167874 79892
rect 167926 79840 167932 79892
rect 167638 79704 167644 79756
rect 167696 79704 167702 79756
rect 167730 79704 167736 79756
rect 167788 79716 167822 79756
rect 167788 79704 167794 79716
rect 167886 79620 167914 79840
rect 167420 79580 167592 79608
rect 167420 79568 167426 79580
rect 167822 79568 167828 79620
rect 167880 79580 167914 79620
rect 167880 79568 167886 79580
rect 166902 79540 166908 79552
rect 166736 79512 166908 79540
rect 166902 79500 166908 79512
rect 166960 79500 166966 79552
rect 166994 79500 167000 79552
rect 167052 79540 167058 79552
rect 167454 79540 167460 79552
rect 167052 79512 167460 79540
rect 167052 79500 167058 79512
rect 167454 79500 167460 79512
rect 167512 79500 167518 79552
rect 166718 79472 166724 79484
rect 166644 79444 166724 79472
rect 165488 79432 165494 79444
rect 166718 79432 166724 79444
rect 166776 79432 166782 79484
rect 167178 79432 167184 79484
rect 167236 79472 167242 79484
rect 167978 79472 168006 79908
rect 168070 79688 168098 79988
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168880 79948 168886 79960
rect 168576 79920 168886 79948
rect 168144 79840 168150 79892
rect 168202 79880 168208 79892
rect 168346 79880 168374 79908
rect 168202 79840 168236 79880
rect 168208 79688 168236 79840
rect 168300 79852 168374 79880
rect 168300 79824 168328 79852
rect 168438 79824 168466 79908
rect 168282 79772 168288 79824
rect 168340 79772 168346 79824
rect 168374 79772 168380 79824
rect 168432 79784 168466 79824
rect 168432 79772 168438 79784
rect 168070 79648 168104 79688
rect 168098 79636 168104 79648
rect 168156 79636 168162 79688
rect 168190 79636 168196 79688
rect 168248 79636 168254 79688
rect 168576 79608 168604 79920
rect 168880 79908 168886 79920
rect 168938 79908 168944 79960
rect 169064 79948 169070 79960
rect 169036 79908 169070 79948
rect 169122 79908 169128 79960
rect 169524 79948 169530 79960
rect 169450 79920 169530 79948
rect 168696 79840 168702 79892
rect 168754 79880 168760 79892
rect 168754 79852 168972 79880
rect 168754 79840 168760 79852
rect 168944 79824 168972 79852
rect 169036 79824 169064 79908
rect 169156 79880 169162 79892
rect 169128 79840 169162 79880
rect 169214 79840 169220 79892
rect 168926 79772 168932 79824
rect 168984 79772 168990 79824
rect 169018 79772 169024 79824
rect 169076 79772 169082 79824
rect 169128 79756 169156 79840
rect 169248 79772 169254 79824
rect 169306 79772 169312 79824
rect 169340 79772 169346 79824
rect 169398 79772 169404 79824
rect 169110 79704 169116 79756
rect 169168 79704 169174 79756
rect 169266 79676 169294 79772
rect 169128 79648 169294 79676
rect 168834 79608 168840 79620
rect 168576 79580 168840 79608
rect 168834 79568 168840 79580
rect 168892 79568 168898 79620
rect 168374 79500 168380 79552
rect 168432 79540 168438 79552
rect 169128 79540 169156 79648
rect 169202 79568 169208 79620
rect 169260 79608 169266 79620
rect 169358 79608 169386 79772
rect 169260 79580 169386 79608
rect 169450 79620 169478 79920
rect 169524 79908 169530 79920
rect 169582 79908 169588 79960
rect 169984 79908 169990 79960
rect 170042 79908 170048 79960
rect 170076 79908 170082 79960
rect 170134 79908 170140 79960
rect 170168 79908 170174 79960
rect 170226 79908 170232 79960
rect 170352 79908 170358 79960
rect 170410 79908 170416 79960
rect 170536 79908 170542 79960
rect 170594 79908 170600 79960
rect 170628 79908 170634 79960
rect 170686 79908 170692 79960
rect 169616 79880 169622 79892
rect 169588 79840 169622 79880
rect 169674 79840 169680 79892
rect 169708 79840 169714 79892
rect 169766 79840 169772 79892
rect 169800 79840 169806 79892
rect 169858 79840 169864 79892
rect 169588 79756 169616 79840
rect 169726 79756 169754 79840
rect 169570 79704 169576 79756
rect 169628 79704 169634 79756
rect 169662 79704 169668 79756
rect 169720 79716 169754 79756
rect 169720 79704 169726 79716
rect 169818 79688 169846 79840
rect 170002 79824 170030 79908
rect 169938 79772 169944 79824
rect 169996 79784 170030 79824
rect 169996 79772 170002 79784
rect 170094 79744 170122 79908
rect 169754 79636 169760 79688
rect 169812 79648 169846 79688
rect 169956 79716 170122 79744
rect 169812 79636 169818 79648
rect 169450 79580 169484 79620
rect 169260 79568 169266 79580
rect 169478 79568 169484 79580
rect 169536 79568 169542 79620
rect 169956 79608 169984 79716
rect 170030 79636 170036 79688
rect 170088 79676 170094 79688
rect 170186 79676 170214 79908
rect 170370 79756 170398 79908
rect 170554 79824 170582 79908
rect 170490 79772 170496 79824
rect 170548 79784 170582 79824
rect 170548 79772 170554 79784
rect 170646 79756 170674 79908
rect 170738 79880 170766 80192
rect 171658 80152 171686 80260
rect 174446 80248 174452 80300
rect 174504 80288 174510 80300
rect 180150 80288 180156 80300
rect 174504 80260 180156 80288
rect 174504 80248 174510 80260
rect 180150 80248 180156 80260
rect 180208 80248 180214 80300
rect 172578 80192 174584 80220
rect 171658 80124 172146 80152
rect 172118 80084 172146 80124
rect 172578 80084 172606 80192
rect 174446 80152 174452 80164
rect 172118 80056 172606 80084
rect 172762 80124 174452 80152
rect 171180 79908 171186 79960
rect 171238 79948 171244 79960
rect 171238 79920 171962 79948
rect 171238 79908 171244 79920
rect 171732 79880 171738 79892
rect 170738 79852 171134 79880
rect 170370 79716 170404 79756
rect 170398 79704 170404 79716
rect 170456 79704 170462 79756
rect 170582 79704 170588 79756
rect 170640 79716 170674 79756
rect 170640 79704 170646 79716
rect 170088 79648 170214 79676
rect 170088 79636 170094 79648
rect 170122 79608 170128 79620
rect 169956 79580 170128 79608
rect 170122 79568 170128 79580
rect 170180 79568 170186 79620
rect 171106 79608 171134 79852
rect 171612 79852 171738 79880
rect 171612 79688 171640 79852
rect 171732 79840 171738 79852
rect 171790 79840 171796 79892
rect 171934 79880 171962 79920
rect 172008 79908 172014 79960
rect 172066 79948 172072 79960
rect 172762 79948 172790 80124
rect 174446 80112 174452 80124
rect 174504 80112 174510 80164
rect 174556 80152 174584 80192
rect 178586 80180 178592 80232
rect 178644 80220 178650 80232
rect 356054 80220 356060 80232
rect 178644 80192 356060 80220
rect 178644 80180 178650 80192
rect 356054 80180 356060 80192
rect 356112 80180 356118 80232
rect 373994 80152 374000 80164
rect 174556 80124 374000 80152
rect 373994 80112 374000 80124
rect 374052 80112 374058 80164
rect 172066 79920 172790 79948
rect 172854 80056 174492 80084
rect 172066 79908 172072 79920
rect 172854 79880 172882 80056
rect 174464 80016 174492 80056
rect 174538 80044 174544 80096
rect 174596 80084 174602 80096
rect 426434 80084 426440 80096
rect 174596 80056 426440 80084
rect 174596 80044 174602 80056
rect 426434 80044 426440 80056
rect 426492 80044 426498 80096
rect 175274 80016 175280 80028
rect 173590 79988 174400 80016
rect 174464 79988 175280 80016
rect 173590 79960 173618 79988
rect 174372 79960 174400 79988
rect 175274 79976 175280 79988
rect 175332 79976 175338 80028
rect 173112 79908 173118 79960
rect 173170 79908 173176 79960
rect 173204 79908 173210 79960
rect 173262 79908 173268 79960
rect 173480 79948 173486 79960
rect 173314 79920 173486 79948
rect 171934 79852 172882 79880
rect 172928 79840 172934 79892
rect 172986 79880 172992 79892
rect 172986 79840 173020 79880
rect 172992 79756 173020 79840
rect 173130 79824 173158 79908
rect 173066 79772 173072 79824
rect 173124 79784 173158 79824
rect 173124 79772 173130 79784
rect 172974 79704 172980 79756
rect 173032 79704 173038 79756
rect 173222 79688 173250 79908
rect 173314 79756 173342 79920
rect 173480 79908 173486 79920
rect 173538 79908 173544 79960
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173756 79908 173762 79960
rect 173814 79908 173820 79960
rect 173848 79908 173854 79960
rect 173906 79948 173912 79960
rect 173906 79908 173940 79948
rect 174032 79908 174038 79960
rect 174090 79908 174096 79960
rect 174354 79908 174360 79960
rect 174412 79908 174418 79960
rect 173388 79840 173394 79892
rect 173446 79880 173452 79892
rect 173774 79880 173802 79908
rect 173446 79852 173572 79880
rect 173774 79852 173848 79880
rect 173446 79840 173452 79852
rect 173544 79756 173572 79852
rect 173314 79716 173348 79756
rect 173342 79704 173348 79716
rect 173400 79704 173406 79756
rect 173526 79704 173532 79756
rect 173584 79704 173590 79756
rect 173820 79744 173848 79852
rect 173912 79824 173940 79908
rect 173894 79772 173900 79824
rect 173952 79772 173958 79824
rect 173820 79716 173940 79744
rect 173912 79688 173940 79716
rect 174050 79688 174078 79908
rect 171594 79636 171600 79688
rect 171652 79636 171658 79688
rect 173158 79636 173164 79688
rect 173216 79648 173250 79688
rect 173216 79636 173222 79648
rect 173894 79636 173900 79688
rect 173952 79636 173958 79688
rect 173986 79636 173992 79688
rect 174044 79648 174078 79688
rect 174044 79636 174050 79648
rect 171502 79608 171508 79620
rect 171106 79580 171508 79608
rect 171502 79568 171508 79580
rect 171560 79568 171566 79620
rect 172054 79568 172060 79620
rect 172112 79608 172118 79620
rect 172514 79608 172520 79620
rect 172112 79580 172520 79608
rect 172112 79568 172118 79580
rect 172514 79568 172520 79580
rect 172572 79568 172578 79620
rect 176286 79608 176292 79620
rect 172624 79580 176292 79608
rect 168432 79512 169156 79540
rect 168432 79500 168438 79512
rect 169846 79500 169852 79552
rect 169904 79540 169910 79552
rect 170306 79540 170312 79552
rect 169904 79512 170312 79540
rect 169904 79500 169910 79512
rect 170306 79500 170312 79512
rect 170364 79500 170370 79552
rect 171594 79500 171600 79552
rect 171652 79540 171658 79552
rect 172624 79540 172652 79580
rect 176286 79568 176292 79580
rect 176344 79568 176350 79620
rect 171652 79512 172652 79540
rect 171652 79500 171658 79512
rect 172698 79500 172704 79552
rect 172756 79540 172762 79552
rect 173066 79540 173072 79552
rect 172756 79512 173072 79540
rect 172756 79500 172762 79512
rect 173066 79500 173072 79512
rect 173124 79500 173130 79552
rect 173710 79500 173716 79552
rect 173768 79540 173774 79552
rect 173768 79512 179414 79540
rect 173768 79500 173774 79512
rect 167236 79444 168006 79472
rect 167236 79432 167242 79444
rect 171318 79432 171324 79484
rect 171376 79472 171382 79484
rect 171376 79444 171732 79472
rect 171376 79432 171382 79444
rect 171704 79404 171732 79444
rect 171778 79432 171784 79484
rect 171836 79472 171842 79484
rect 177022 79472 177028 79484
rect 171836 79444 177028 79472
rect 171836 79432 171842 79444
rect 177022 79432 177028 79444
rect 177080 79432 177086 79484
rect 179386 79472 179414 79512
rect 179386 79444 180794 79472
rect 180242 79404 180248 79416
rect 143592 79376 161152 79404
rect 161216 79376 171640 79404
rect 171704 79376 180248 79404
rect 143592 79364 143598 79376
rect 152550 79336 152556 79348
rect 136284 79308 152556 79336
rect 128780 79296 128786 79308
rect 152550 79296 152556 79308
rect 152608 79296 152614 79348
rect 153102 79296 153108 79348
rect 153160 79336 153166 79348
rect 160738 79336 160744 79348
rect 153160 79308 160744 79336
rect 153160 79296 153166 79308
rect 160738 79296 160744 79308
rect 160796 79296 160802 79348
rect 161124 79336 161152 79376
rect 171134 79336 171140 79348
rect 161124 79308 171140 79336
rect 171134 79296 171140 79308
rect 171192 79296 171198 79348
rect 171612 79336 171640 79376
rect 180242 79364 180248 79376
rect 180300 79364 180306 79416
rect 180766 79404 180794 79444
rect 527174 79404 527180 79416
rect 180766 79376 527180 79404
rect 527174 79364 527180 79376
rect 527232 79364 527238 79416
rect 171962 79336 171968 79348
rect 171612 79308 171968 79336
rect 171962 79296 171968 79308
rect 172020 79296 172026 79348
rect 172514 79296 172520 79348
rect 172572 79336 172578 79348
rect 580074 79336 580080 79348
rect 172572 79308 580080 79336
rect 172572 79296 172578 79308
rect 580074 79296 580080 79308
rect 580132 79296 580138 79348
rect 120626 79228 120632 79280
rect 120684 79268 120690 79280
rect 166994 79268 167000 79280
rect 120684 79240 167000 79268
rect 120684 79228 120690 79240
rect 166994 79228 167000 79240
rect 167052 79228 167058 79280
rect 168006 79228 168012 79280
rect 168064 79268 168070 79280
rect 173894 79268 173900 79280
rect 168064 79240 173900 79268
rect 168064 79228 168070 79240
rect 173894 79228 173900 79240
rect 173952 79228 173958 79280
rect 143534 79200 143540 79212
rect 120552 79172 130148 79200
rect 128722 79132 128728 79144
rect 116636 79104 118694 79132
rect 120460 79104 128728 79132
rect 116636 79092 116642 79104
rect 118666 78996 118694 79104
rect 128722 79092 128728 79104
rect 128780 79092 128786 79144
rect 130120 79132 130148 79172
rect 135226 79172 143540 79200
rect 135226 79132 135254 79172
rect 143534 79160 143540 79172
rect 143592 79160 143598 79212
rect 153194 79160 153200 79212
rect 153252 79200 153258 79212
rect 157702 79200 157708 79212
rect 153252 79172 157708 79200
rect 153252 79160 153258 79172
rect 157702 79160 157708 79172
rect 157760 79160 157766 79212
rect 160370 79160 160376 79212
rect 160428 79200 160434 79212
rect 160554 79200 160560 79212
rect 160428 79172 160560 79200
rect 160428 79160 160434 79172
rect 160554 79160 160560 79172
rect 160612 79160 160618 79212
rect 160738 79160 160744 79212
rect 160796 79200 160802 79212
rect 171318 79200 171324 79212
rect 160796 79172 171324 79200
rect 160796 79160 160802 79172
rect 171318 79160 171324 79172
rect 171376 79160 171382 79212
rect 173986 79200 173992 79212
rect 171520 79172 173992 79200
rect 171520 79132 171548 79172
rect 173986 79160 173992 79172
rect 174044 79160 174050 79212
rect 172330 79132 172336 79144
rect 130120 79104 135254 79132
rect 137986 79104 171548 79132
rect 171612 79104 172336 79132
rect 127894 79024 127900 79076
rect 127952 79064 127958 79076
rect 137094 79064 137100 79076
rect 127952 79036 137100 79064
rect 127952 79024 127958 79036
rect 137094 79024 137100 79036
rect 137152 79024 137158 79076
rect 137986 78996 138014 79104
rect 152642 79024 152648 79076
rect 152700 79064 152706 79076
rect 153010 79064 153016 79076
rect 152700 79036 153016 79064
rect 152700 79024 152706 79036
rect 153010 79024 153016 79036
rect 153068 79024 153074 79076
rect 154574 79024 154580 79076
rect 154632 79064 154638 79076
rect 171612 79064 171640 79104
rect 172330 79092 172336 79104
rect 172388 79092 172394 79144
rect 172422 79092 172428 79144
rect 172480 79132 172486 79144
rect 175918 79132 175924 79144
rect 172480 79104 175924 79132
rect 172480 79092 172486 79104
rect 175918 79092 175924 79104
rect 175976 79092 175982 79144
rect 154632 79036 171640 79064
rect 154632 79024 154638 79036
rect 171686 79024 171692 79076
rect 171744 79064 171750 79076
rect 398190 79064 398196 79076
rect 171744 79036 398196 79064
rect 171744 79024 171750 79036
rect 398190 79024 398196 79036
rect 398248 79024 398254 79076
rect 118666 78968 138014 78996
rect 159174 78956 159180 79008
rect 159232 78996 159238 79008
rect 430574 78996 430580 79008
rect 159232 78968 430580 78996
rect 159232 78956 159238 78968
rect 430574 78956 430580 78968
rect 430632 78956 430638 79008
rect 127434 78888 127440 78940
rect 127492 78928 127498 78940
rect 127710 78928 127716 78940
rect 127492 78900 127716 78928
rect 127492 78888 127498 78900
rect 127710 78888 127716 78900
rect 127768 78888 127774 78940
rect 137094 78888 137100 78940
rect 137152 78928 137158 78940
rect 148318 78928 148324 78940
rect 137152 78900 148324 78928
rect 137152 78888 137158 78900
rect 148318 78888 148324 78900
rect 148376 78888 148382 78940
rect 151906 78888 151912 78940
rect 151964 78928 151970 78940
rect 152642 78928 152648 78940
rect 151964 78900 152648 78928
rect 151964 78888 151970 78900
rect 152642 78888 152648 78900
rect 152700 78888 152706 78940
rect 157794 78888 157800 78940
rect 157852 78928 157858 78940
rect 164050 78928 164056 78940
rect 157852 78900 164056 78928
rect 157852 78888 157858 78900
rect 164050 78888 164056 78900
rect 164108 78888 164114 78940
rect 171410 78928 171416 78940
rect 164942 78900 171416 78928
rect 125962 78820 125968 78872
rect 126020 78860 126026 78872
rect 127526 78860 127532 78872
rect 126020 78832 127532 78860
rect 126020 78820 126026 78832
rect 127526 78820 127532 78832
rect 127584 78820 127590 78872
rect 152550 78820 152556 78872
rect 152608 78860 152614 78872
rect 163130 78860 163136 78872
rect 152608 78832 163136 78860
rect 152608 78820 152614 78832
rect 163130 78820 163136 78832
rect 163188 78820 163194 78872
rect 127710 78752 127716 78804
rect 127768 78792 127774 78804
rect 129366 78792 129372 78804
rect 127768 78764 129372 78792
rect 127768 78752 127774 78764
rect 129366 78752 129372 78764
rect 129424 78752 129430 78804
rect 152090 78752 152096 78804
rect 152148 78792 152154 78804
rect 154390 78792 154396 78804
rect 152148 78764 154396 78792
rect 152148 78752 152154 78764
rect 154390 78752 154396 78764
rect 154448 78752 154454 78804
rect 154942 78752 154948 78804
rect 155000 78792 155006 78804
rect 155126 78792 155132 78804
rect 155000 78764 155132 78792
rect 155000 78752 155006 78764
rect 155126 78752 155132 78764
rect 155184 78752 155190 78804
rect 156414 78752 156420 78804
rect 156472 78792 156478 78804
rect 160370 78792 160376 78804
rect 156472 78764 160376 78792
rect 156472 78752 156478 78764
rect 160370 78752 160376 78764
rect 160428 78752 160434 78804
rect 161566 78752 161572 78804
rect 161624 78792 161630 78804
rect 164942 78792 164970 78900
rect 171410 78888 171416 78900
rect 171468 78888 171474 78940
rect 172054 78888 172060 78940
rect 172112 78928 172118 78940
rect 173250 78928 173256 78940
rect 172112 78900 173256 78928
rect 172112 78888 172118 78900
rect 173250 78888 173256 78900
rect 173308 78888 173314 78940
rect 176102 78888 176108 78940
rect 176160 78928 176166 78940
rect 504358 78928 504364 78940
rect 176160 78900 504364 78928
rect 176160 78888 176166 78900
rect 504358 78888 504364 78900
rect 504416 78888 504422 78940
rect 165706 78820 165712 78872
rect 165764 78860 165770 78872
rect 166166 78860 166172 78872
rect 165764 78832 166172 78860
rect 165764 78820 165770 78832
rect 166166 78820 166172 78832
rect 166224 78820 166230 78872
rect 167454 78820 167460 78872
rect 167512 78860 167518 78872
rect 532694 78860 532700 78872
rect 167512 78832 532700 78860
rect 167512 78820 167518 78832
rect 532694 78820 532700 78832
rect 532752 78820 532758 78872
rect 161624 78764 164970 78792
rect 161624 78752 161630 78764
rect 168466 78752 168472 78804
rect 168524 78792 168530 78804
rect 168650 78792 168656 78804
rect 168524 78764 168656 78792
rect 168524 78752 168530 78764
rect 168650 78752 168656 78764
rect 168708 78752 168714 78804
rect 168926 78752 168932 78804
rect 168984 78792 168990 78804
rect 554774 78792 554780 78804
rect 168984 78764 554780 78792
rect 168984 78752 168990 78764
rect 554774 78752 554780 78764
rect 554832 78752 554838 78804
rect 151446 78684 151452 78736
rect 151504 78724 151510 78736
rect 153194 78724 153200 78736
rect 151504 78696 153200 78724
rect 151504 78684 151510 78696
rect 153194 78684 153200 78696
rect 153252 78684 153258 78736
rect 164234 78684 164240 78736
rect 164292 78724 164298 78736
rect 169570 78724 169576 78736
rect 164292 78696 169576 78724
rect 164292 78684 164298 78696
rect 169570 78684 169576 78696
rect 169628 78684 169634 78736
rect 170306 78684 170312 78736
rect 170364 78724 170370 78736
rect 557534 78724 557540 78736
rect 170364 78696 557540 78724
rect 170364 78684 170370 78696
rect 557534 78684 557540 78696
rect 557592 78684 557598 78736
rect 128354 78616 128360 78668
rect 128412 78656 128418 78668
rect 131574 78656 131580 78668
rect 128412 78628 131580 78656
rect 128412 78616 128418 78628
rect 131574 78616 131580 78628
rect 131632 78616 131638 78668
rect 135530 78616 135536 78668
rect 135588 78656 135594 78668
rect 135898 78656 135904 78668
rect 135588 78628 135904 78656
rect 135588 78616 135594 78628
rect 135898 78616 135904 78628
rect 135956 78616 135962 78668
rect 136818 78616 136824 78668
rect 136876 78656 136882 78668
rect 137370 78656 137376 78668
rect 136876 78628 137376 78656
rect 136876 78616 136882 78628
rect 137370 78616 137376 78628
rect 137428 78616 137434 78668
rect 138106 78616 138112 78668
rect 138164 78656 138170 78668
rect 138566 78656 138572 78668
rect 138164 78628 138572 78656
rect 138164 78616 138170 78628
rect 138566 78616 138572 78628
rect 138624 78616 138630 78668
rect 140866 78616 140872 78668
rect 140924 78656 140930 78668
rect 141510 78656 141516 78668
rect 140924 78628 141516 78656
rect 140924 78616 140930 78628
rect 141510 78616 141516 78628
rect 141568 78616 141574 78668
rect 153378 78616 153384 78668
rect 153436 78656 153442 78668
rect 153654 78656 153660 78668
rect 153436 78628 153660 78656
rect 153436 78616 153442 78628
rect 153654 78616 153660 78628
rect 153712 78616 153718 78668
rect 160922 78616 160928 78668
rect 160980 78656 160986 78668
rect 162394 78656 162400 78668
rect 160980 78628 162400 78656
rect 160980 78616 160986 78628
rect 162394 78616 162400 78628
rect 162452 78616 162458 78668
rect 164418 78616 164424 78668
rect 164476 78656 164482 78668
rect 164602 78656 164608 78668
rect 164476 78628 164608 78656
rect 164476 78616 164482 78628
rect 164602 78616 164608 78628
rect 164660 78616 164666 78668
rect 398098 78656 398104 78668
rect 190426 78628 398104 78656
rect 128538 78588 128544 78600
rect 124186 78560 128544 78588
rect 122190 78412 122196 78464
rect 122248 78452 122254 78464
rect 124186 78452 124214 78560
rect 128538 78548 128544 78560
rect 128596 78548 128602 78600
rect 137002 78548 137008 78600
rect 137060 78588 137066 78600
rect 137186 78588 137192 78600
rect 137060 78560 137192 78588
rect 137060 78548 137066 78560
rect 137186 78548 137192 78560
rect 137244 78548 137250 78600
rect 138934 78548 138940 78600
rect 138992 78588 138998 78600
rect 139118 78588 139124 78600
rect 138992 78560 139124 78588
rect 138992 78548 138998 78560
rect 139118 78548 139124 78560
rect 139176 78548 139182 78600
rect 150434 78548 150440 78600
rect 150492 78588 150498 78600
rect 156966 78588 156972 78600
rect 150492 78560 156972 78588
rect 150492 78548 150498 78560
rect 156966 78548 156972 78560
rect 157024 78548 157030 78600
rect 159634 78548 159640 78600
rect 159692 78588 159698 78600
rect 168006 78588 168012 78600
rect 159692 78560 168012 78588
rect 159692 78548 159698 78560
rect 168006 78548 168012 78560
rect 168064 78548 168070 78600
rect 174170 78588 174176 78600
rect 168116 78560 174176 78588
rect 164602 78520 164608 78532
rect 159100 78492 164608 78520
rect 122248 78424 124214 78452
rect 122248 78412 122254 78424
rect 128538 78412 128544 78464
rect 128596 78452 128602 78464
rect 132862 78452 132868 78464
rect 128596 78424 132868 78452
rect 128596 78412 128602 78424
rect 132862 78412 132868 78424
rect 132920 78412 132926 78464
rect 147674 78412 147680 78464
rect 147732 78452 147738 78464
rect 159100 78452 159128 78492
rect 164602 78480 164608 78492
rect 164660 78480 164666 78532
rect 166166 78480 166172 78532
rect 166224 78520 166230 78532
rect 166350 78520 166356 78532
rect 166224 78492 166356 78520
rect 166224 78480 166230 78492
rect 166350 78480 166356 78492
rect 166408 78480 166414 78532
rect 166994 78480 167000 78532
rect 167052 78520 167058 78532
rect 168116 78520 168144 78560
rect 174170 78548 174176 78560
rect 174228 78548 174234 78600
rect 175642 78548 175648 78600
rect 175700 78588 175706 78600
rect 190426 78588 190454 78628
rect 398098 78616 398104 78628
rect 398156 78616 398162 78668
rect 175700 78560 190454 78588
rect 175700 78548 175706 78560
rect 167052 78492 168144 78520
rect 167052 78480 167058 78492
rect 172146 78480 172152 78532
rect 172204 78520 172210 78532
rect 180058 78520 180064 78532
rect 172204 78492 180064 78520
rect 172204 78480 172210 78492
rect 180058 78480 180064 78492
rect 180116 78480 180122 78532
rect 397546 78520 397552 78532
rect 183526 78492 397552 78520
rect 147732 78424 159128 78452
rect 147732 78412 147738 78424
rect 160370 78412 160376 78464
rect 160428 78452 160434 78464
rect 172054 78452 172060 78464
rect 160428 78424 172060 78452
rect 160428 78412 160434 78424
rect 172054 78412 172060 78424
rect 172112 78412 172118 78464
rect 173250 78412 173256 78464
rect 173308 78452 173314 78464
rect 183526 78452 183554 78492
rect 397546 78480 397552 78492
rect 397604 78480 397610 78532
rect 173308 78424 183554 78452
rect 173308 78412 173314 78424
rect 116578 78344 116584 78396
rect 116636 78384 116642 78396
rect 129182 78384 129188 78396
rect 116636 78356 129188 78384
rect 116636 78344 116642 78356
rect 129182 78344 129188 78356
rect 129240 78344 129246 78396
rect 141050 78344 141056 78396
rect 141108 78384 141114 78396
rect 171594 78384 171600 78396
rect 141108 78356 171600 78384
rect 141108 78344 141114 78356
rect 171594 78344 171600 78356
rect 171652 78344 171658 78396
rect 171870 78344 171876 78396
rect 171928 78384 171934 78396
rect 179966 78384 179972 78396
rect 171928 78356 179972 78384
rect 171928 78344 171934 78356
rect 179966 78344 179972 78356
rect 180024 78344 180030 78396
rect 114554 78276 114560 78328
rect 114612 78316 114618 78328
rect 134426 78316 134432 78328
rect 114612 78288 134432 78316
rect 114612 78276 114618 78288
rect 134426 78276 134432 78288
rect 134484 78276 134490 78328
rect 138382 78276 138388 78328
rect 138440 78316 138446 78328
rect 138750 78316 138756 78328
rect 138440 78288 138756 78316
rect 138440 78276 138446 78288
rect 138750 78276 138756 78288
rect 138808 78276 138814 78328
rect 139946 78276 139952 78328
rect 140004 78316 140010 78328
rect 178034 78316 178040 78328
rect 140004 78288 178040 78316
rect 140004 78276 140010 78288
rect 178034 78276 178040 78288
rect 178092 78276 178098 78328
rect 113818 78208 113824 78260
rect 113876 78248 113882 78260
rect 125318 78248 125324 78260
rect 113876 78220 125324 78248
rect 113876 78208 113882 78220
rect 125318 78208 125324 78220
rect 125376 78208 125382 78260
rect 131574 78208 131580 78260
rect 131632 78248 131638 78260
rect 132126 78248 132132 78260
rect 131632 78220 132132 78248
rect 131632 78208 131638 78220
rect 132126 78208 132132 78220
rect 132184 78208 132190 78260
rect 134058 78208 134064 78260
rect 134116 78248 134122 78260
rect 134242 78248 134248 78260
rect 134116 78220 134248 78248
rect 134116 78208 134122 78220
rect 134242 78208 134248 78220
rect 134300 78208 134306 78260
rect 141050 78208 141056 78260
rect 141108 78248 141114 78260
rect 141602 78248 141608 78260
rect 141108 78220 141608 78248
rect 141108 78208 141114 78220
rect 141602 78208 141608 78220
rect 141660 78208 141666 78260
rect 161566 78208 161572 78260
rect 161624 78248 161630 78260
rect 162118 78248 162124 78260
rect 161624 78220 162124 78248
rect 161624 78208 161630 78220
rect 162118 78208 162124 78220
rect 162176 78208 162182 78260
rect 162394 78208 162400 78260
rect 162452 78248 162458 78260
rect 242158 78248 242164 78260
rect 162452 78220 242164 78248
rect 162452 78208 162458 78220
rect 242158 78208 242164 78220
rect 242216 78208 242222 78260
rect 110414 78140 110420 78192
rect 110472 78180 110478 78192
rect 122926 78180 122932 78192
rect 110472 78152 122932 78180
rect 110472 78140 110478 78152
rect 122926 78140 122932 78152
rect 122984 78140 122990 78192
rect 123294 78140 123300 78192
rect 123352 78180 123358 78192
rect 123352 78152 124214 78180
rect 123352 78140 123358 78152
rect 107654 78072 107660 78124
rect 107712 78112 107718 78124
rect 123386 78112 123392 78124
rect 107712 78084 123392 78112
rect 107712 78072 107718 78084
rect 123386 78072 123392 78084
rect 123444 78072 123450 78124
rect 124186 78112 124214 78152
rect 126054 78140 126060 78192
rect 126112 78180 126118 78192
rect 126330 78180 126336 78192
rect 126112 78152 126336 78180
rect 126112 78140 126118 78152
rect 126330 78140 126336 78152
rect 126388 78140 126394 78192
rect 126422 78140 126428 78192
rect 126480 78180 126486 78192
rect 130470 78180 130476 78192
rect 126480 78152 130476 78180
rect 126480 78140 126486 78152
rect 130470 78140 130476 78152
rect 130528 78140 130534 78192
rect 133874 78140 133880 78192
rect 133932 78180 133938 78192
rect 135990 78180 135996 78192
rect 133932 78152 135996 78180
rect 133932 78140 133938 78152
rect 135990 78140 135996 78152
rect 136048 78140 136054 78192
rect 144178 78140 144184 78192
rect 144236 78180 144242 78192
rect 152550 78180 152556 78192
rect 144236 78152 152556 78180
rect 144236 78140 144242 78152
rect 152550 78140 152556 78152
rect 152608 78140 152614 78192
rect 159358 78140 159364 78192
rect 159416 78180 159422 78192
rect 162946 78180 162952 78192
rect 159416 78152 162952 78180
rect 159416 78140 159422 78152
rect 162946 78140 162952 78152
rect 163004 78140 163010 78192
rect 304258 78180 304264 78192
rect 163056 78152 304264 78180
rect 124186 78084 127388 78112
rect 93118 78004 93124 78056
rect 93176 78044 93182 78056
rect 125962 78044 125968 78056
rect 93176 78016 125968 78044
rect 93176 78004 93182 78016
rect 125962 78004 125968 78016
rect 126020 78004 126026 78056
rect 127360 78044 127388 78084
rect 127894 78072 127900 78124
rect 127952 78112 127958 78124
rect 135438 78112 135444 78124
rect 127952 78084 135444 78112
rect 127952 78072 127958 78084
rect 135438 78072 135444 78084
rect 135496 78072 135502 78124
rect 160922 78112 160928 78124
rect 152476 78084 160928 78112
rect 132770 78044 132776 78056
rect 127360 78016 132776 78044
rect 132770 78004 132776 78016
rect 132828 78004 132834 78056
rect 134242 78004 134248 78056
rect 134300 78044 134306 78056
rect 134886 78044 134892 78056
rect 134300 78016 134892 78044
rect 134300 78004 134306 78016
rect 134886 78004 134892 78016
rect 134944 78004 134950 78056
rect 135990 78004 135996 78056
rect 136048 78044 136054 78056
rect 136174 78044 136180 78056
rect 136048 78016 136180 78044
rect 136048 78004 136054 78016
rect 136174 78004 136180 78016
rect 136232 78004 136238 78056
rect 89714 77936 89720 77988
rect 89772 77976 89778 77988
rect 123294 77976 123300 77988
rect 89772 77948 123300 77976
rect 89772 77936 89778 77948
rect 123294 77936 123300 77948
rect 123352 77936 123358 77988
rect 124950 77936 124956 77988
rect 125008 77976 125014 77988
rect 127066 77976 127072 77988
rect 125008 77948 127072 77976
rect 125008 77936 125014 77948
rect 127066 77936 127072 77948
rect 127124 77936 127130 77988
rect 127434 77936 127440 77988
rect 127492 77976 127498 77988
rect 127618 77976 127624 77988
rect 127492 77948 127624 77976
rect 127492 77936 127498 77948
rect 127618 77936 127624 77948
rect 127676 77936 127682 77988
rect 130194 77936 130200 77988
rect 130252 77976 130258 77988
rect 130378 77976 130384 77988
rect 130252 77948 130384 77976
rect 130252 77936 130258 77948
rect 130378 77936 130384 77948
rect 130436 77936 130442 77988
rect 131298 77936 131304 77988
rect 131356 77976 131362 77988
rect 132034 77976 132040 77988
rect 131356 77948 132040 77976
rect 131356 77936 131362 77948
rect 132034 77936 132040 77948
rect 132092 77936 132098 77988
rect 134426 77936 134432 77988
rect 134484 77976 134490 77988
rect 134794 77976 134800 77988
rect 134484 77948 134800 77976
rect 134484 77936 134490 77948
rect 134794 77936 134800 77948
rect 134852 77936 134858 77988
rect 139670 77936 139676 77988
rect 139728 77976 139734 77988
rect 152476 77976 152504 78084
rect 160922 78072 160928 78084
rect 160980 78072 160986 78124
rect 161658 78072 161664 78124
rect 161716 78112 161722 78124
rect 163056 78112 163084 78152
rect 304258 78140 304264 78152
rect 304316 78140 304322 78192
rect 161716 78084 163084 78112
rect 164206 78084 169524 78112
rect 161716 78072 161722 78084
rect 157058 78004 157064 78056
rect 157116 78044 157122 78056
rect 164206 78044 164234 78084
rect 157116 78016 164234 78044
rect 157116 78004 157122 78016
rect 139728 77948 152504 77976
rect 139728 77936 139734 77948
rect 155494 77936 155500 77988
rect 155552 77976 155558 77988
rect 159634 77976 159640 77988
rect 155552 77948 159640 77976
rect 155552 77936 155558 77948
rect 159634 77936 159640 77948
rect 159692 77936 159698 77988
rect 162946 77936 162952 77988
rect 163004 77976 163010 77988
rect 169386 77976 169392 77988
rect 163004 77948 169392 77976
rect 163004 77936 163010 77948
rect 169386 77936 169392 77948
rect 169444 77936 169450 77988
rect 125318 77868 125324 77920
rect 125376 77908 125382 77920
rect 133414 77908 133420 77920
rect 125376 77880 133420 77908
rect 125376 77868 125382 77880
rect 133414 77868 133420 77880
rect 133472 77868 133478 77920
rect 142062 77868 142068 77920
rect 142120 77908 142126 77920
rect 152182 77908 152188 77920
rect 142120 77880 152188 77908
rect 142120 77868 142126 77880
rect 152182 77868 152188 77880
rect 152240 77868 152246 77920
rect 164234 77908 164240 77920
rect 152292 77880 164240 77908
rect 120074 77800 120080 77852
rect 120132 77840 120138 77852
rect 124030 77840 124036 77852
rect 120132 77812 124036 77840
rect 120132 77800 120138 77812
rect 124030 77800 124036 77812
rect 124088 77800 124094 77852
rect 124122 77800 124128 77852
rect 124180 77840 124186 77852
rect 135346 77840 135352 77852
rect 124180 77812 135352 77840
rect 124180 77800 124186 77812
rect 135346 77800 135352 77812
rect 135404 77800 135410 77852
rect 144914 77800 144920 77852
rect 144972 77840 144978 77852
rect 152292 77840 152320 77880
rect 164234 77868 164240 77880
rect 164292 77868 164298 77920
rect 169496 77908 169524 78084
rect 169570 78072 169576 78124
rect 169628 78112 169634 78124
rect 498194 78112 498200 78124
rect 169628 78084 498200 78112
rect 169628 78072 169634 78084
rect 498194 78072 498200 78084
rect 498252 78072 498258 78124
rect 170582 78004 170588 78056
rect 170640 78044 170646 78056
rect 574738 78044 574744 78056
rect 170640 78016 574744 78044
rect 170640 78004 170646 78016
rect 574738 78004 574744 78016
rect 574796 78004 574802 78056
rect 170766 77936 170772 77988
rect 170824 77976 170830 77988
rect 581086 77976 581092 77988
rect 170824 77948 581092 77976
rect 170824 77936 170830 77948
rect 581086 77936 581092 77948
rect 581144 77936 581150 77988
rect 171962 77908 171968 77920
rect 169496 77880 171968 77908
rect 171962 77868 171968 77880
rect 172020 77868 172026 77920
rect 172054 77868 172060 77920
rect 172112 77908 172118 77920
rect 173618 77908 173624 77920
rect 172112 77880 173624 77908
rect 172112 77868 172118 77880
rect 173618 77868 173624 77880
rect 173676 77868 173682 77920
rect 173986 77868 173992 77920
rect 174044 77908 174050 77920
rect 174446 77908 174452 77920
rect 174044 77880 174452 77908
rect 174044 77868 174050 77880
rect 174446 77868 174452 77880
rect 174504 77868 174510 77920
rect 144972 77812 152320 77840
rect 144972 77800 144978 77812
rect 152550 77800 152556 77852
rect 152608 77840 152614 77852
rect 162118 77840 162124 77852
rect 152608 77812 162124 77840
rect 152608 77800 152614 77812
rect 162118 77800 162124 77812
rect 162176 77800 162182 77852
rect 165890 77800 165896 77852
rect 165948 77840 165954 77852
rect 170582 77840 170588 77852
rect 165948 77812 170588 77840
rect 165948 77800 165954 77812
rect 170582 77800 170588 77812
rect 170640 77800 170646 77852
rect 171318 77800 171324 77852
rect 171376 77840 171382 77852
rect 172422 77840 172428 77852
rect 171376 77812 172428 77840
rect 171376 77800 171382 77812
rect 172422 77800 172428 77812
rect 172480 77800 172486 77852
rect 129182 77732 129188 77784
rect 129240 77772 129246 77784
rect 129826 77772 129832 77784
rect 129240 77744 129832 77772
rect 129240 77732 129246 77744
rect 129826 77732 129832 77744
rect 129884 77732 129890 77784
rect 131298 77732 131304 77784
rect 131356 77772 131362 77784
rect 131758 77772 131764 77784
rect 131356 77744 131764 77772
rect 131356 77732 131362 77744
rect 131758 77732 131764 77744
rect 131816 77732 131822 77784
rect 159174 77732 159180 77784
rect 159232 77772 159238 77784
rect 159232 77744 162716 77772
rect 159232 77732 159238 77744
rect 158898 77664 158904 77716
rect 158956 77704 158962 77716
rect 162688 77704 162716 77744
rect 164050 77732 164056 77784
rect 164108 77772 164114 77784
rect 172238 77772 172244 77784
rect 164108 77744 172244 77772
rect 164108 77732 164114 77744
rect 172238 77732 172244 77744
rect 172296 77732 172302 77784
rect 171778 77704 171784 77716
rect 158956 77676 162624 77704
rect 162688 77676 171784 77704
rect 158956 77664 158962 77676
rect 125134 77596 125140 77648
rect 125192 77636 125198 77648
rect 126698 77636 126704 77648
rect 125192 77608 126704 77636
rect 125192 77596 125198 77608
rect 126698 77596 126704 77608
rect 126756 77596 126762 77648
rect 155862 77596 155868 77648
rect 155920 77636 155926 77648
rect 162486 77636 162492 77648
rect 155920 77608 162492 77636
rect 155920 77596 155926 77608
rect 162486 77596 162492 77608
rect 162544 77596 162550 77648
rect 162596 77636 162624 77676
rect 171778 77664 171784 77676
rect 171836 77664 171842 77716
rect 171686 77636 171692 77648
rect 162596 77608 171692 77636
rect 171686 77596 171692 77608
rect 171744 77596 171750 77648
rect 123386 77528 123392 77580
rect 123444 77568 123450 77580
rect 129734 77568 129740 77580
rect 123444 77540 129740 77568
rect 123444 77528 123450 77540
rect 129734 77528 129740 77540
rect 129792 77528 129798 77580
rect 147674 77528 147680 77580
rect 147732 77568 147738 77580
rect 148042 77568 148048 77580
rect 147732 77540 148048 77568
rect 147732 77528 147738 77540
rect 148042 77528 148048 77540
rect 148100 77528 148106 77580
rect 154666 77528 154672 77580
rect 154724 77568 154730 77580
rect 158254 77568 158260 77580
rect 154724 77540 158260 77568
rect 154724 77528 154730 77540
rect 158254 77528 158260 77540
rect 158312 77528 158318 77580
rect 159910 77528 159916 77580
rect 159968 77568 159974 77580
rect 172054 77568 172060 77580
rect 159968 77540 172060 77568
rect 159968 77528 159974 77540
rect 172054 77528 172060 77540
rect 172112 77528 172118 77580
rect 122926 77460 122932 77512
rect 122984 77500 122990 77512
rect 134058 77500 134064 77512
rect 122984 77472 134064 77500
rect 122984 77460 122990 77472
rect 134058 77460 134064 77472
rect 134116 77460 134122 77512
rect 152182 77460 152188 77512
rect 152240 77500 152246 77512
rect 152826 77500 152832 77512
rect 152240 77472 152832 77500
rect 152240 77460 152246 77472
rect 152826 77460 152832 77472
rect 152884 77460 152890 77512
rect 154482 77460 154488 77512
rect 154540 77500 154546 77512
rect 158622 77500 158628 77512
rect 154540 77472 158628 77500
rect 154540 77460 154546 77472
rect 158622 77460 158628 77472
rect 158680 77460 158686 77512
rect 163130 77460 163136 77512
rect 163188 77500 163194 77512
rect 173342 77500 173348 77512
rect 163188 77472 173348 77500
rect 163188 77460 163194 77472
rect 173342 77460 173348 77472
rect 173400 77460 173406 77512
rect 123570 77392 123576 77444
rect 123628 77432 123634 77444
rect 134978 77432 134984 77444
rect 123628 77404 134984 77432
rect 123628 77392 123634 77404
rect 134978 77392 134984 77404
rect 135036 77392 135042 77444
rect 154022 77392 154028 77444
rect 154080 77432 154086 77444
rect 154080 77404 154574 77432
rect 154080 77392 154086 77404
rect 120810 77324 120816 77376
rect 120868 77364 120874 77376
rect 128078 77364 128084 77376
rect 120868 77336 128084 77364
rect 120868 77324 120874 77336
rect 128078 77324 128084 77336
rect 128136 77324 128142 77376
rect 150342 77324 150348 77376
rect 150400 77364 150406 77376
rect 153102 77364 153108 77376
rect 150400 77336 153108 77364
rect 150400 77324 150406 77336
rect 153102 77324 153108 77336
rect 153160 77324 153166 77376
rect 153378 77324 153384 77376
rect 153436 77364 153442 77376
rect 154114 77364 154120 77376
rect 153436 77336 154120 77364
rect 153436 77324 153442 77336
rect 154114 77324 154120 77336
rect 154172 77324 154178 77376
rect 154546 77364 154574 77404
rect 154666 77392 154672 77444
rect 154724 77432 154730 77444
rect 155310 77432 155316 77444
rect 154724 77404 155316 77432
rect 154724 77392 154730 77404
rect 155310 77392 155316 77404
rect 155368 77392 155374 77444
rect 157426 77392 157432 77444
rect 157484 77432 157490 77444
rect 157978 77432 157984 77444
rect 157484 77404 157984 77432
rect 157484 77392 157490 77404
rect 157978 77392 157984 77404
rect 158036 77392 158042 77444
rect 169386 77392 169392 77444
rect 169444 77432 169450 77444
rect 175918 77432 175924 77444
rect 169444 77404 175924 77432
rect 169444 77392 169450 77404
rect 175918 77392 175924 77404
rect 175976 77392 175982 77444
rect 180058 77392 180064 77444
rect 180116 77432 180122 77444
rect 396718 77432 396724 77444
rect 180116 77404 396724 77432
rect 180116 77392 180122 77404
rect 396718 77392 396724 77404
rect 396776 77392 396782 77444
rect 155218 77364 155224 77376
rect 154546 77336 155224 77364
rect 155218 77324 155224 77336
rect 155276 77324 155282 77376
rect 155402 77324 155408 77376
rect 155460 77364 155466 77376
rect 155678 77364 155684 77376
rect 155460 77336 155684 77364
rect 155460 77324 155466 77336
rect 155678 77324 155684 77336
rect 155736 77324 155742 77376
rect 127066 77256 127072 77308
rect 127124 77296 127130 77308
rect 127894 77296 127900 77308
rect 127124 77268 127900 77296
rect 127124 77256 127130 77268
rect 127894 77256 127900 77268
rect 127952 77256 127958 77308
rect 130470 77256 130476 77308
rect 130528 77296 130534 77308
rect 135806 77296 135812 77308
rect 130528 77268 135812 77296
rect 130528 77256 130534 77268
rect 135806 77256 135812 77268
rect 135864 77256 135870 77308
rect 149514 77256 149520 77308
rect 149572 77296 149578 77308
rect 149698 77296 149704 77308
rect 149572 77268 149704 77296
rect 149572 77256 149578 77268
rect 149698 77256 149704 77268
rect 149756 77256 149762 77308
rect 152182 77256 152188 77308
rect 152240 77296 152246 77308
rect 152458 77296 152464 77308
rect 152240 77268 152464 77296
rect 152240 77256 152246 77268
rect 152458 77256 152464 77268
rect 152516 77256 152522 77308
rect 154206 77256 154212 77308
rect 154264 77296 154270 77308
rect 155494 77296 155500 77308
rect 154264 77268 155500 77296
rect 154264 77256 154270 77268
rect 155494 77256 155500 77268
rect 155552 77256 155558 77308
rect 156414 77256 156420 77308
rect 156472 77296 156478 77308
rect 156690 77296 156696 77308
rect 156472 77268 156696 77296
rect 156472 77256 156478 77268
rect 156690 77256 156696 77268
rect 156748 77256 156754 77308
rect 119430 77188 119436 77240
rect 119488 77228 119494 77240
rect 172882 77228 172888 77240
rect 119488 77200 172888 77228
rect 119488 77188 119494 77200
rect 172882 77188 172888 77200
rect 172940 77188 172946 77240
rect 143166 77120 143172 77172
rect 143224 77160 143230 77172
rect 226334 77160 226340 77172
rect 143224 77132 226340 77160
rect 143224 77120 143230 77132
rect 226334 77120 226340 77132
rect 226392 77120 226398 77172
rect 168834 77092 168840 77104
rect 152384 77064 168840 77092
rect 123478 76984 123484 77036
rect 123536 77024 123542 77036
rect 132310 77024 132316 77036
rect 123536 76996 132316 77024
rect 123536 76984 123542 76996
rect 132310 76984 132316 76996
rect 132368 76984 132374 77036
rect 147950 76984 147956 77036
rect 148008 77024 148014 77036
rect 148410 77024 148416 77036
rect 148008 76996 148416 77024
rect 148008 76984 148014 76996
rect 148410 76984 148416 76996
rect 148468 76984 148474 77036
rect 149238 76984 149244 77036
rect 149296 77024 149302 77036
rect 149974 77024 149980 77036
rect 149296 76996 149980 77024
rect 149296 76984 149302 76996
rect 149974 76984 149980 76996
rect 150032 76984 150038 77036
rect 124858 76916 124864 76968
rect 124916 76956 124922 76968
rect 135162 76956 135168 76968
rect 124916 76928 135168 76956
rect 124916 76916 124922 76928
rect 135162 76916 135168 76928
rect 135220 76916 135226 76968
rect 149146 76916 149152 76968
rect 149204 76956 149210 76968
rect 149606 76956 149612 76968
rect 149204 76928 149612 76956
rect 149204 76916 149210 76928
rect 149606 76916 149612 76928
rect 149664 76916 149670 76968
rect 150158 76916 150164 76968
rect 150216 76956 150222 76968
rect 152384 76956 152412 77064
rect 168834 77052 168840 77064
rect 168892 77052 168898 77104
rect 171778 77052 171784 77104
rect 171836 77092 171842 77104
rect 249794 77092 249800 77104
rect 171836 77064 249800 77092
rect 171836 77052 171842 77064
rect 249794 77052 249800 77064
rect 249852 77052 249858 77104
rect 247034 77024 247040 77036
rect 150216 76928 152412 76956
rect 152476 76996 164234 77024
rect 150216 76916 150222 76928
rect 118694 76848 118700 76900
rect 118752 76888 118758 76900
rect 134610 76888 134616 76900
rect 118752 76860 134616 76888
rect 118752 76848 118758 76860
rect 134610 76848 134616 76860
rect 134668 76848 134674 76900
rect 144822 76848 144828 76900
rect 144880 76888 144886 76900
rect 152476 76888 152504 76996
rect 164206 76956 164234 76996
rect 167104 76996 247040 77024
rect 167104 76956 167132 76996
rect 247034 76984 247040 76996
rect 247092 76984 247098 77036
rect 164206 76928 167132 76956
rect 168834 76916 168840 76968
rect 168892 76956 168898 76968
rect 260834 76956 260840 76968
rect 168892 76928 260840 76956
rect 168892 76916 168898 76928
rect 260834 76916 260840 76928
rect 260892 76916 260898 76968
rect 144880 76860 152504 76888
rect 144880 76848 144886 76860
rect 164602 76848 164608 76900
rect 164660 76888 164666 76900
rect 284294 76888 284300 76900
rect 164660 76860 284300 76888
rect 164660 76848 164666 76860
rect 284294 76848 284300 76860
rect 284352 76848 284358 76900
rect 102134 76780 102140 76832
rect 102192 76820 102198 76832
rect 132678 76820 132684 76832
rect 102192 76792 132684 76820
rect 102192 76780 102198 76792
rect 132678 76780 132684 76792
rect 132736 76780 132742 76832
rect 143718 76780 143724 76832
rect 143776 76820 143782 76832
rect 144362 76820 144368 76832
rect 143776 76792 144368 76820
rect 143776 76780 143782 76792
rect 144362 76780 144368 76792
rect 144420 76780 144426 76832
rect 148594 76780 148600 76832
rect 148652 76820 148658 76832
rect 296714 76820 296720 76832
rect 148652 76792 296720 76820
rect 148652 76780 148658 76792
rect 296714 76780 296720 76792
rect 296772 76780 296778 76832
rect 70394 76712 70400 76764
rect 70452 76752 70458 76764
rect 131206 76752 131212 76764
rect 70452 76724 131212 76752
rect 70452 76712 70458 76724
rect 131206 76712 131212 76724
rect 131264 76712 131270 76764
rect 135162 76712 135168 76764
rect 135220 76752 135226 76764
rect 138014 76752 138020 76764
rect 135220 76724 138020 76752
rect 135220 76712 135226 76724
rect 138014 76712 138020 76724
rect 138072 76712 138078 76764
rect 148042 76712 148048 76764
rect 148100 76752 148106 76764
rect 148318 76752 148324 76764
rect 148100 76724 148324 76752
rect 148100 76712 148106 76724
rect 148318 76712 148324 76724
rect 148376 76712 148382 76764
rect 149238 76712 149244 76764
rect 149296 76752 149302 76764
rect 149882 76752 149888 76764
rect 149296 76724 149888 76752
rect 149296 76712 149302 76724
rect 149882 76712 149888 76724
rect 149940 76712 149946 76764
rect 152274 76712 152280 76764
rect 152332 76752 152338 76764
rect 152734 76752 152740 76764
rect 152332 76724 152740 76752
rect 152332 76712 152338 76724
rect 152734 76712 152740 76724
rect 152792 76712 152798 76764
rect 157610 76712 157616 76764
rect 157668 76752 157674 76764
rect 157886 76752 157892 76764
rect 157668 76724 157892 76752
rect 157668 76712 157674 76724
rect 157886 76712 157892 76724
rect 157944 76712 157950 76764
rect 164234 76712 164240 76764
rect 164292 76752 164298 76764
rect 171778 76752 171784 76764
rect 164292 76724 171784 76752
rect 164292 76712 164298 76724
rect 171778 76712 171784 76724
rect 171836 76712 171842 76764
rect 172330 76712 172336 76764
rect 172388 76752 172394 76764
rect 376754 76752 376760 76764
rect 172388 76724 376760 76752
rect 172388 76712 172394 76724
rect 376754 76712 376760 76724
rect 376812 76712 376818 76764
rect 93854 76644 93860 76696
rect 93912 76684 93918 76696
rect 128538 76684 128544 76696
rect 93912 76656 128544 76684
rect 93912 76644 93918 76656
rect 128538 76644 128544 76656
rect 128596 76644 128602 76696
rect 137922 76644 137928 76696
rect 137980 76684 137986 76696
rect 144362 76684 144368 76696
rect 137980 76656 144368 76684
rect 137980 76644 137986 76656
rect 144362 76644 144368 76656
rect 144420 76644 144426 76696
rect 147858 76644 147864 76696
rect 147916 76684 147922 76696
rect 148226 76684 148232 76696
rect 147916 76656 148232 76684
rect 147916 76644 147922 76656
rect 148226 76644 148232 76656
rect 148284 76644 148290 76696
rect 154850 76644 154856 76696
rect 154908 76684 154914 76696
rect 375374 76684 375380 76696
rect 154908 76656 375380 76684
rect 154908 76644 154914 76656
rect 375374 76644 375380 76656
rect 375432 76644 375438 76696
rect 69014 76576 69020 76628
rect 69072 76616 69078 76628
rect 130930 76616 130936 76628
rect 69072 76588 130936 76616
rect 69072 76576 69078 76588
rect 130930 76576 130936 76588
rect 130988 76576 130994 76628
rect 157610 76576 157616 76628
rect 157668 76616 157674 76628
rect 158070 76616 158076 76628
rect 157668 76588 158076 76616
rect 157668 76576 157674 76588
rect 158070 76576 158076 76588
rect 158128 76576 158134 76628
rect 160094 76576 160100 76628
rect 160152 76616 160158 76628
rect 444374 76616 444380 76628
rect 160152 76588 444380 76616
rect 160152 76576 160158 76588
rect 444374 76576 444380 76588
rect 444432 76576 444438 76628
rect 6914 76508 6920 76560
rect 6972 76548 6978 76560
rect 124766 76548 124772 76560
rect 6972 76520 124772 76548
rect 6972 76508 6978 76520
rect 124766 76508 124772 76520
rect 124824 76508 124830 76560
rect 147674 76508 147680 76560
rect 147732 76548 147738 76560
rect 147858 76548 147864 76560
rect 147732 76520 147864 76548
rect 147732 76508 147738 76520
rect 147858 76508 147864 76520
rect 147916 76508 147922 76560
rect 154850 76508 154856 76560
rect 154908 76548 154914 76560
rect 155402 76548 155408 76560
rect 154908 76520 155408 76548
rect 154908 76508 154914 76520
rect 155402 76508 155408 76520
rect 155460 76508 155466 76560
rect 165614 76508 165620 76560
rect 165672 76548 165678 76560
rect 170674 76548 170680 76560
rect 165672 76520 170680 76548
rect 165672 76508 165678 76520
rect 170674 76508 170680 76520
rect 170732 76508 170738 76560
rect 171594 76508 171600 76560
rect 171652 76548 171658 76560
rect 171870 76548 171876 76560
rect 171652 76520 171876 76548
rect 171652 76508 171658 76520
rect 171870 76508 171876 76520
rect 171928 76508 171934 76560
rect 558914 76548 558920 76560
rect 172486 76520 558920 76548
rect 132954 76440 132960 76492
rect 133012 76480 133018 76492
rect 133230 76480 133236 76492
rect 133012 76452 133236 76480
rect 133012 76440 133018 76452
rect 133230 76440 133236 76452
rect 133288 76440 133294 76492
rect 140406 76440 140412 76492
rect 140464 76480 140470 76492
rect 140464 76452 157334 76480
rect 140464 76440 140470 76452
rect 147674 76372 147680 76424
rect 147732 76412 147738 76424
rect 148502 76412 148508 76424
rect 147732 76384 148508 76412
rect 147732 76372 147738 76384
rect 148502 76372 148508 76384
rect 148560 76372 148566 76424
rect 139302 76304 139308 76356
rect 139360 76344 139366 76356
rect 140406 76344 140412 76356
rect 139360 76316 140412 76344
rect 139360 76304 139366 76316
rect 140406 76304 140412 76316
rect 140464 76304 140470 76356
rect 147030 76236 147036 76288
rect 147088 76236 147094 76288
rect 157306 76276 157334 76452
rect 168558 76440 168564 76492
rect 168616 76480 168622 76492
rect 168926 76480 168932 76492
rect 168616 76452 168932 76480
rect 168616 76440 168622 76452
rect 168926 76440 168932 76452
rect 168984 76440 168990 76492
rect 169018 76440 169024 76492
rect 169076 76480 169082 76492
rect 172486 76480 172514 76520
rect 558914 76508 558920 76520
rect 558972 76508 558978 76560
rect 190454 76480 190460 76492
rect 169076 76452 172514 76480
rect 176626 76452 190460 76480
rect 169076 76440 169082 76452
rect 170950 76372 170956 76424
rect 171008 76412 171014 76424
rect 173342 76412 173348 76424
rect 171008 76384 173348 76412
rect 171008 76372 171014 76384
rect 173342 76372 173348 76384
rect 173400 76372 173406 76424
rect 171410 76304 171416 76356
rect 171468 76344 171474 76356
rect 172330 76344 172336 76356
rect 171468 76316 172336 76344
rect 171468 76304 171474 76316
rect 172330 76304 172336 76316
rect 172388 76304 172394 76356
rect 176626 76276 176654 76452
rect 190454 76440 190460 76452
rect 190512 76440 190518 76492
rect 157306 76248 176654 76276
rect 146846 76208 146852 76220
rect 146404 76180 146852 76208
rect 140774 76032 140780 76084
rect 140832 76072 140838 76084
rect 141142 76072 141148 76084
rect 140832 76044 141148 76072
rect 140832 76032 140838 76044
rect 141142 76032 141148 76044
rect 141200 76032 141206 76084
rect 145006 76032 145012 76084
rect 145064 76072 145070 76084
rect 145064 76044 145144 76072
rect 145064 76032 145070 76044
rect 145116 76016 145144 76044
rect 124030 75964 124036 76016
rect 124088 76004 124094 76016
rect 124088 75976 124260 76004
rect 124088 75964 124094 75976
rect 120718 75896 120724 75948
rect 120776 75936 120782 75948
rect 120776 75908 124168 75936
rect 120776 75896 120782 75908
rect 124140 75800 124168 75908
rect 124232 75868 124260 75976
rect 145098 75964 145104 76016
rect 145156 75964 145162 76016
rect 145374 75964 145380 76016
rect 145432 76004 145438 76016
rect 145650 76004 145656 76016
rect 145432 75976 145656 76004
rect 145432 75964 145438 75976
rect 145650 75964 145656 75976
rect 145708 75964 145714 76016
rect 139670 75896 139676 75948
rect 139728 75936 139734 75948
rect 140038 75936 140044 75948
rect 139728 75908 140044 75936
rect 139728 75896 139734 75908
rect 140038 75896 140044 75908
rect 140096 75896 140102 75948
rect 141142 75896 141148 75948
rect 141200 75936 141206 75948
rect 141694 75936 141700 75948
rect 141200 75908 141700 75936
rect 141200 75896 141206 75908
rect 141694 75896 141700 75908
rect 141752 75896 141758 75948
rect 144178 75896 144184 75948
rect 144236 75936 144242 75948
rect 144730 75936 144736 75948
rect 144236 75908 144736 75936
rect 144236 75896 144242 75908
rect 144730 75896 144736 75908
rect 144788 75896 144794 75948
rect 146404 75936 146432 76180
rect 146846 76168 146852 76180
rect 146904 76168 146910 76220
rect 147048 76208 147076 76236
rect 147048 76180 147168 76208
rect 146662 76100 146668 76152
rect 146720 76140 146726 76152
rect 147030 76140 147036 76152
rect 146720 76112 147036 76140
rect 146720 76100 146726 76112
rect 147030 76100 147036 76112
rect 147088 76100 147094 76152
rect 146478 76032 146484 76084
rect 146536 76072 146542 76084
rect 146846 76072 146852 76084
rect 146536 76044 146852 76072
rect 146536 76032 146542 76044
rect 146846 76032 146852 76044
rect 146904 76032 146910 76084
rect 146662 75964 146668 76016
rect 146720 76004 146726 76016
rect 147140 76004 147168 76180
rect 160094 76168 160100 76220
rect 160152 76208 160158 76220
rect 160554 76208 160560 76220
rect 160152 76180 160560 76208
rect 160152 76168 160158 76180
rect 160554 76168 160560 76180
rect 160612 76168 160618 76220
rect 165798 76168 165804 76220
rect 165856 76208 165862 76220
rect 166810 76208 166816 76220
rect 165856 76180 166816 76208
rect 165856 76168 165862 76180
rect 166810 76168 166816 76180
rect 166868 76168 166874 76220
rect 160646 76140 160652 76152
rect 160480 76112 160652 76140
rect 146720 75976 147168 76004
rect 146720 75964 146726 75976
rect 150434 75964 150440 76016
rect 150492 76004 150498 76016
rect 150618 76004 150624 76016
rect 150492 75976 150624 76004
rect 150492 75964 150498 75976
rect 150618 75964 150624 75976
rect 150676 75964 150682 76016
rect 146478 75936 146484 75948
rect 146404 75908 146484 75936
rect 146478 75896 146484 75908
rect 146536 75896 146542 75948
rect 146570 75896 146576 75948
rect 146628 75936 146634 75948
rect 147214 75936 147220 75948
rect 146628 75908 147220 75936
rect 146628 75896 146634 75908
rect 147214 75896 147220 75908
rect 147272 75896 147278 75948
rect 158898 75896 158904 75948
rect 158956 75936 158962 75948
rect 159450 75936 159456 75948
rect 158956 75908 159456 75936
rect 158956 75896 158962 75908
rect 159450 75896 159456 75908
rect 159508 75896 159514 75948
rect 160480 75936 160508 76112
rect 160646 76100 160652 76112
rect 160704 76100 160710 76152
rect 161750 76100 161756 76152
rect 161808 76140 161814 76152
rect 161934 76140 161940 76152
rect 161808 76112 161940 76140
rect 161808 76100 161814 76112
rect 161934 76100 161940 76112
rect 161992 76100 161998 76152
rect 163406 76140 163412 76152
rect 162872 76112 163412 76140
rect 162872 76084 162900 76112
rect 163406 76100 163412 76112
rect 163464 76100 163470 76152
rect 162854 76032 162860 76084
rect 162912 76032 162918 76084
rect 162946 76032 162952 76084
rect 163004 76072 163010 76084
rect 163958 76072 163964 76084
rect 163004 76044 163964 76072
rect 163004 76032 163010 76044
rect 163958 76032 163964 76044
rect 164016 76032 164022 76084
rect 161750 75964 161756 76016
rect 161808 76004 161814 76016
rect 162026 76004 162032 76016
rect 161808 75976 162032 76004
rect 161808 75964 161814 75976
rect 162026 75964 162032 75976
rect 162084 75964 162090 76016
rect 163130 75964 163136 76016
rect 163188 76004 163194 76016
rect 163866 76004 163872 76016
rect 163188 75976 163872 76004
rect 163188 75964 163194 75976
rect 163866 75964 163872 75976
rect 163924 75964 163930 76016
rect 160554 75936 160560 75948
rect 160480 75908 160560 75936
rect 160554 75896 160560 75908
rect 160612 75896 160618 75948
rect 161474 75896 161480 75948
rect 161532 75936 161538 75948
rect 162210 75936 162216 75948
rect 161532 75908 162216 75936
rect 161532 75896 161538 75908
rect 162210 75896 162216 75908
rect 162268 75896 162274 75948
rect 163406 75896 163412 75948
rect 163464 75936 163470 75948
rect 163682 75936 163688 75948
rect 163464 75908 163688 75936
rect 163464 75896 163470 75908
rect 163682 75896 163688 75908
rect 163740 75896 163746 75948
rect 164602 75896 164608 75948
rect 164660 75936 164666 75948
rect 165246 75936 165252 75948
rect 164660 75908 165252 75936
rect 164660 75896 164666 75908
rect 165246 75896 165252 75908
rect 165304 75896 165310 75948
rect 165430 75896 165436 75948
rect 165488 75936 165494 75948
rect 165798 75936 165804 75948
rect 165488 75908 165804 75936
rect 165488 75896 165494 75908
rect 165798 75896 165804 75908
rect 165856 75896 165862 75948
rect 165890 75896 165896 75948
rect 165948 75936 165954 75948
rect 166626 75936 166632 75948
rect 165948 75908 166632 75936
rect 165948 75896 165954 75908
rect 166626 75896 166632 75908
rect 166684 75896 166690 75948
rect 166902 75896 166908 75948
rect 166960 75936 166966 75948
rect 167362 75936 167368 75948
rect 166960 75908 167368 75936
rect 166960 75896 166966 75908
rect 167362 75896 167368 75908
rect 167420 75896 167426 75948
rect 167454 75896 167460 75948
rect 167512 75936 167518 75948
rect 167730 75936 167736 75948
rect 167512 75908 167736 75936
rect 167512 75896 167518 75908
rect 167730 75896 167736 75908
rect 167788 75896 167794 75948
rect 172698 75868 172704 75880
rect 124232 75840 172704 75868
rect 172698 75828 172704 75840
rect 172756 75828 172762 75880
rect 172514 75800 172520 75812
rect 124140 75772 172520 75800
rect 172514 75760 172520 75772
rect 172572 75760 172578 75812
rect 139946 75692 139952 75744
rect 140004 75732 140010 75744
rect 140222 75732 140228 75744
rect 140004 75704 140228 75732
rect 140004 75692 140010 75704
rect 140222 75692 140228 75704
rect 140280 75692 140286 75744
rect 159082 75692 159088 75744
rect 159140 75732 159146 75744
rect 159818 75732 159824 75744
rect 159140 75704 159824 75732
rect 159140 75692 159146 75704
rect 159818 75692 159824 75704
rect 159876 75692 159882 75744
rect 160094 75692 160100 75744
rect 160152 75732 160158 75744
rect 161014 75732 161020 75744
rect 160152 75704 161020 75732
rect 160152 75692 160158 75704
rect 161014 75692 161020 75704
rect 161072 75692 161078 75744
rect 167362 75692 167368 75744
rect 167420 75732 167426 75744
rect 167638 75732 167644 75744
rect 167420 75704 167644 75732
rect 167420 75692 167426 75704
rect 167638 75692 167644 75704
rect 167696 75692 167702 75744
rect 139578 75624 139584 75676
rect 139636 75664 139642 75676
rect 140130 75664 140136 75676
rect 139636 75636 140136 75664
rect 139636 75624 139642 75636
rect 140130 75624 140136 75636
rect 140188 75624 140194 75676
rect 157334 75624 157340 75676
rect 157392 75664 157398 75676
rect 158162 75664 158168 75676
rect 157392 75636 158168 75664
rect 157392 75624 157398 75636
rect 158162 75624 158168 75636
rect 158220 75624 158226 75676
rect 132034 75596 132040 75608
rect 118666 75568 132040 75596
rect 75914 75420 75920 75472
rect 75972 75460 75978 75472
rect 118666 75460 118694 75568
rect 132034 75556 132040 75568
rect 132092 75556 132098 75608
rect 121454 75488 121460 75540
rect 121512 75528 121518 75540
rect 134610 75528 134616 75540
rect 121512 75500 134616 75528
rect 121512 75488 121518 75500
rect 134610 75488 134616 75500
rect 134668 75488 134674 75540
rect 162578 75488 162584 75540
rect 162636 75528 162642 75540
rect 162636 75500 168374 75528
rect 162636 75488 162642 75500
rect 75972 75432 118694 75460
rect 75972 75420 75978 75432
rect 127158 75420 127164 75472
rect 127216 75460 127222 75472
rect 127710 75460 127716 75472
rect 127216 75432 127716 75460
rect 127216 75420 127222 75432
rect 127710 75420 127716 75432
rect 127768 75420 127774 75472
rect 159726 75420 159732 75472
rect 159784 75460 159790 75472
rect 168346 75460 168374 75500
rect 169938 75488 169944 75540
rect 169996 75528 170002 75540
rect 170306 75528 170312 75540
rect 169996 75500 170312 75528
rect 169996 75488 170002 75500
rect 170306 75488 170312 75500
rect 170364 75488 170370 75540
rect 431954 75460 431960 75472
rect 159784 75432 164050 75460
rect 168346 75432 431960 75460
rect 159784 75420 159790 75432
rect 51074 75352 51080 75404
rect 51132 75392 51138 75404
rect 128998 75392 129004 75404
rect 51132 75364 129004 75392
rect 51132 75352 51138 75364
rect 128998 75352 129004 75364
rect 129056 75352 129062 75404
rect 137094 75352 137100 75404
rect 137152 75392 137158 75404
rect 137738 75392 137744 75404
rect 137152 75364 137744 75392
rect 137152 75352 137158 75364
rect 137738 75352 137744 75364
rect 137796 75352 137802 75404
rect 150802 75352 150808 75404
rect 150860 75392 150866 75404
rect 163774 75392 163780 75404
rect 150860 75364 163780 75392
rect 150860 75352 150866 75364
rect 163774 75352 163780 75364
rect 163832 75352 163838 75404
rect 164022 75392 164050 75432
rect 431954 75420 431960 75432
rect 432012 75420 432018 75472
rect 438854 75392 438860 75404
rect 164022 75364 438860 75392
rect 438854 75352 438860 75364
rect 438912 75352 438918 75404
rect 49694 75284 49700 75336
rect 49752 75324 49758 75336
rect 127158 75324 127164 75336
rect 49752 75296 127164 75324
rect 49752 75284 49758 75296
rect 127158 75284 127164 75296
rect 127216 75284 127222 75336
rect 127250 75284 127256 75336
rect 127308 75324 127314 75336
rect 128078 75324 128084 75336
rect 127308 75296 128084 75324
rect 127308 75284 127314 75296
rect 128078 75284 128084 75296
rect 128136 75284 128142 75336
rect 128538 75284 128544 75336
rect 128596 75324 128602 75336
rect 129642 75324 129648 75336
rect 128596 75296 129648 75324
rect 128596 75284 128602 75296
rect 129642 75284 129648 75296
rect 129700 75284 129706 75336
rect 132678 75284 132684 75336
rect 132736 75324 132742 75336
rect 133598 75324 133604 75336
rect 132736 75296 133604 75324
rect 132736 75284 132742 75296
rect 133598 75284 133604 75296
rect 133656 75284 133662 75336
rect 135346 75284 135352 75336
rect 135404 75324 135410 75336
rect 135622 75324 135628 75336
rect 135404 75296 135628 75324
rect 135404 75284 135410 75296
rect 135622 75284 135628 75296
rect 135680 75284 135686 75336
rect 135806 75284 135812 75336
rect 135864 75324 135870 75336
rect 136450 75324 136456 75336
rect 135864 75296 136456 75324
rect 135864 75284 135870 75296
rect 136450 75284 136456 75296
rect 136508 75284 136514 75336
rect 164878 75284 164884 75336
rect 164936 75324 164942 75336
rect 481634 75324 481640 75336
rect 164936 75296 481640 75324
rect 164936 75284 164942 75296
rect 481634 75284 481640 75296
rect 481692 75284 481698 75336
rect 46934 75216 46940 75268
rect 46992 75256 46998 75268
rect 46992 75228 128354 75256
rect 46992 75216 46998 75228
rect 26234 75148 26240 75200
rect 26292 75188 26298 75200
rect 26292 75160 118694 75188
rect 26292 75148 26298 75160
rect 118666 75052 118694 75160
rect 125962 75148 125968 75200
rect 126020 75188 126026 75200
rect 126882 75188 126888 75200
rect 126020 75160 126888 75188
rect 126020 75148 126026 75160
rect 126882 75148 126888 75160
rect 126940 75148 126946 75200
rect 127158 75148 127164 75200
rect 127216 75188 127222 75200
rect 127802 75188 127808 75200
rect 127216 75160 127808 75188
rect 127216 75148 127222 75160
rect 127802 75148 127808 75160
rect 127860 75148 127866 75200
rect 127066 75080 127072 75132
rect 127124 75120 127130 75132
rect 127434 75120 127440 75132
rect 127124 75092 127440 75120
rect 127124 75080 127130 75092
rect 127434 75080 127440 75092
rect 127492 75080 127498 75132
rect 128326 75120 128354 75228
rect 128722 75216 128728 75268
rect 128780 75256 128786 75268
rect 129090 75256 129096 75268
rect 128780 75228 129096 75256
rect 128780 75216 128786 75228
rect 129090 75216 129096 75228
rect 129148 75216 129154 75268
rect 130010 75216 130016 75268
rect 130068 75256 130074 75268
rect 130654 75256 130660 75268
rect 130068 75228 130660 75256
rect 130068 75216 130074 75228
rect 130654 75216 130660 75228
rect 130712 75216 130718 75268
rect 131390 75216 131396 75268
rect 131448 75256 131454 75268
rect 131942 75256 131948 75268
rect 131448 75228 131948 75256
rect 131448 75216 131454 75228
rect 131942 75216 131948 75228
rect 132000 75216 132006 75268
rect 133046 75216 133052 75268
rect 133104 75256 133110 75268
rect 133782 75256 133788 75268
rect 133104 75228 133788 75256
rect 133104 75216 133110 75228
rect 133782 75216 133788 75228
rect 133840 75216 133846 75268
rect 134150 75216 134156 75268
rect 134208 75256 134214 75268
rect 134518 75256 134524 75268
rect 134208 75228 134524 75256
rect 134208 75216 134214 75228
rect 134518 75216 134524 75228
rect 134576 75216 134582 75268
rect 135714 75216 135720 75268
rect 135772 75256 135778 75268
rect 136266 75256 136272 75268
rect 135772 75228 136272 75256
rect 135772 75216 135778 75228
rect 136266 75216 136272 75228
rect 136324 75216 136330 75268
rect 137094 75216 137100 75268
rect 137152 75256 137158 75268
rect 137462 75256 137468 75268
rect 137152 75228 137468 75256
rect 137152 75216 137158 75228
rect 137462 75216 137468 75228
rect 137520 75216 137526 75268
rect 138290 75216 138296 75268
rect 138348 75256 138354 75268
rect 138474 75256 138480 75268
rect 138348 75228 138480 75256
rect 138348 75216 138354 75228
rect 138474 75216 138480 75228
rect 138532 75216 138538 75268
rect 150802 75216 150808 75268
rect 150860 75256 150866 75268
rect 151170 75256 151176 75268
rect 150860 75228 151176 75256
rect 150860 75216 150866 75228
rect 151170 75216 151176 75228
rect 151228 75216 151234 75268
rect 153194 75216 153200 75268
rect 153252 75256 153258 75268
rect 154114 75256 154120 75268
rect 153252 75228 154120 75256
rect 153252 75216 153258 75228
rect 154114 75216 154120 75228
rect 154172 75216 154178 75268
rect 163866 75216 163872 75268
rect 163924 75256 163930 75268
rect 489914 75256 489920 75268
rect 163924 75228 489920 75256
rect 163924 75216 163930 75228
rect 489914 75216 489920 75228
rect 489972 75216 489978 75268
rect 128630 75148 128636 75200
rect 128688 75188 128694 75200
rect 129550 75188 129556 75200
rect 128688 75160 129556 75188
rect 128688 75148 128694 75160
rect 129550 75148 129556 75160
rect 129608 75148 129614 75200
rect 129734 75148 129740 75200
rect 129792 75188 129798 75200
rect 130470 75188 130476 75200
rect 129792 75160 130476 75188
rect 129792 75148 129798 75160
rect 130470 75148 130476 75160
rect 130528 75148 130534 75200
rect 131206 75148 131212 75200
rect 131264 75188 131270 75200
rect 132126 75188 132132 75200
rect 131264 75160 132132 75188
rect 131264 75148 131270 75160
rect 132126 75148 132132 75160
rect 132184 75148 132190 75200
rect 132770 75148 132776 75200
rect 132828 75188 132834 75200
rect 133690 75188 133696 75200
rect 132828 75160 133696 75188
rect 132828 75148 132834 75160
rect 133690 75148 133696 75160
rect 133748 75148 133754 75200
rect 135622 75148 135628 75200
rect 135680 75188 135686 75200
rect 135990 75188 135996 75200
rect 135680 75160 135996 75188
rect 135680 75148 135686 75160
rect 135990 75148 135996 75160
rect 136048 75148 136054 75200
rect 150618 75148 150624 75200
rect 150676 75188 150682 75200
rect 151078 75188 151084 75200
rect 150676 75160 151084 75188
rect 150676 75148 150682 75160
rect 151078 75148 151084 75160
rect 151136 75148 151142 75200
rect 156230 75148 156236 75200
rect 156288 75188 156294 75200
rect 156506 75188 156512 75200
rect 156288 75160 156512 75188
rect 156288 75148 156294 75160
rect 156506 75148 156512 75160
rect 156564 75148 156570 75200
rect 169754 75148 169760 75200
rect 169812 75188 169818 75200
rect 170030 75188 170036 75200
rect 169812 75160 170036 75188
rect 169812 75148 169818 75160
rect 170030 75148 170036 75160
rect 170088 75148 170094 75200
rect 564434 75188 564440 75200
rect 176626 75160 564440 75188
rect 129366 75120 129372 75132
rect 128326 75092 129372 75120
rect 129366 75080 129372 75092
rect 129424 75080 129430 75132
rect 135438 75080 135444 75132
rect 135496 75120 135502 75132
rect 136358 75120 136364 75132
rect 135496 75092 136364 75120
rect 135496 75080 135502 75092
rect 136358 75080 136364 75092
rect 136416 75080 136422 75132
rect 138290 75080 138296 75132
rect 138348 75120 138354 75132
rect 138566 75120 138572 75132
rect 138348 75092 138572 75120
rect 138348 75080 138354 75092
rect 138566 75080 138572 75092
rect 138624 75080 138630 75132
rect 151906 75080 151912 75132
rect 151964 75120 151970 75132
rect 152458 75120 152464 75132
rect 151964 75092 152464 75120
rect 151964 75080 151970 75092
rect 152458 75080 152464 75092
rect 152516 75080 152522 75132
rect 168834 75080 168840 75132
rect 168892 75120 168898 75132
rect 169202 75120 169208 75132
rect 168892 75092 169208 75120
rect 168892 75080 168898 75092
rect 169202 75080 169208 75092
rect 169260 75080 169266 75132
rect 127986 75052 127992 75064
rect 118666 75024 127992 75052
rect 127986 75012 127992 75024
rect 128044 75012 128050 75064
rect 156046 75012 156052 75064
rect 156104 75052 156110 75064
rect 156506 75052 156512 75064
rect 156104 75024 156512 75052
rect 156104 75012 156110 75024
rect 156506 75012 156512 75024
rect 156564 75012 156570 75064
rect 169754 75012 169760 75064
rect 169812 75052 169818 75064
rect 170214 75052 170220 75064
rect 169812 75024 170220 75052
rect 169812 75012 169818 75024
rect 170214 75012 170220 75024
rect 170272 75012 170278 75064
rect 127434 74944 127440 74996
rect 127492 74984 127498 74996
rect 128262 74984 128268 74996
rect 127492 74956 128268 74984
rect 127492 74944 127498 74956
rect 128262 74944 128268 74956
rect 128320 74944 128326 74996
rect 151906 74944 151912 74996
rect 151964 74984 151970 74996
rect 153010 74984 153016 74996
rect 151964 74956 153016 74984
rect 151964 74944 151970 74956
rect 153010 74944 153016 74956
rect 153068 74944 153074 74996
rect 158806 74944 158812 74996
rect 158864 74984 158870 74996
rect 159266 74984 159272 74996
rect 158864 74956 159272 74984
rect 158864 74944 158870 74956
rect 159266 74944 159272 74956
rect 159324 74944 159330 74996
rect 169294 74944 169300 74996
rect 169352 74984 169358 74996
rect 176626 74984 176654 75160
rect 564434 75148 564440 75160
rect 564492 75148 564498 75200
rect 169352 74956 176654 74984
rect 169352 74944 169358 74956
rect 156046 74876 156052 74928
rect 156104 74916 156110 74928
rect 156782 74916 156788 74928
rect 156104 74888 156788 74916
rect 156104 74876 156110 74888
rect 156782 74876 156788 74888
rect 156840 74876 156846 74928
rect 130470 74468 130476 74520
rect 130528 74508 130534 74520
rect 135254 74508 135260 74520
rect 130528 74480 135260 74508
rect 130528 74468 130534 74480
rect 135254 74468 135260 74480
rect 135312 74468 135318 74520
rect 138750 74468 138756 74520
rect 138808 74508 138814 74520
rect 140130 74508 140136 74520
rect 138808 74480 140136 74508
rect 138808 74468 138814 74480
rect 140130 74468 140136 74480
rect 140188 74468 140194 74520
rect 142246 74128 142252 74180
rect 142304 74168 142310 74180
rect 142798 74168 142804 74180
rect 142304 74140 142804 74168
rect 142304 74128 142310 74140
rect 142798 74128 142804 74140
rect 142856 74128 142862 74180
rect 4154 73992 4160 74044
rect 4212 74032 4218 74044
rect 126330 74032 126336 74044
rect 4212 74004 126336 74032
rect 4212 73992 4218 74004
rect 126330 73992 126336 74004
rect 126388 73992 126394 74044
rect 118786 73924 118792 73976
rect 118844 73964 118850 73976
rect 134426 73964 134432 73976
rect 118844 73936 134432 73964
rect 118844 73924 118850 73936
rect 134426 73924 134432 73936
rect 134484 73924 134490 73976
rect 141878 73924 141884 73976
rect 141936 73964 141942 73976
rect 209774 73964 209780 73976
rect 141936 73936 209780 73964
rect 141936 73924 141942 73936
rect 209774 73924 209780 73936
rect 209832 73924 209838 73976
rect 60734 73856 60740 73908
rect 60792 73896 60798 73908
rect 130194 73896 130200 73908
rect 60792 73868 130200 73896
rect 60792 73856 60798 73868
rect 130194 73856 130200 73868
rect 130252 73856 130258 73908
rect 147306 73856 147312 73908
rect 147364 73896 147370 73908
rect 223574 73896 223580 73908
rect 147364 73868 223580 73896
rect 147364 73856 147370 73868
rect 223574 73856 223580 73868
rect 223632 73856 223638 73908
rect 153194 73788 153200 73840
rect 153252 73828 153258 73840
rect 318794 73828 318800 73840
rect 153252 73800 318800 73828
rect 153252 73788 153258 73800
rect 318794 73788 318800 73800
rect 318852 73788 318858 73840
rect 145006 73720 145012 73772
rect 145064 73760 145070 73772
rect 145834 73760 145840 73772
rect 145064 73732 145840 73760
rect 145064 73720 145070 73732
rect 145834 73720 145840 73732
rect 145892 73720 145898 73772
rect 137554 73516 137560 73568
rect 137612 73556 137618 73568
rect 142982 73556 142988 73568
rect 137612 73528 142988 73556
rect 137612 73516 137618 73528
rect 142982 73516 142988 73528
rect 143040 73516 143046 73568
rect 161658 73448 161664 73500
rect 161716 73488 161722 73500
rect 162302 73488 162308 73500
rect 161716 73460 162308 73488
rect 161716 73448 161722 73460
rect 162302 73448 162308 73460
rect 162360 73448 162366 73500
rect 126238 73176 126244 73228
rect 126296 73216 126302 73228
rect 130838 73216 130844 73228
rect 126296 73188 130844 73216
rect 126296 73176 126302 73188
rect 130838 73176 130844 73188
rect 130896 73176 130902 73228
rect 171042 73108 171048 73160
rect 171100 73148 171106 73160
rect 580166 73148 580172 73160
rect 171100 73120 580172 73148
rect 171100 73108 171106 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 145466 72904 145472 72956
rect 145524 72944 145530 72956
rect 145926 72944 145932 72956
rect 145524 72916 145932 72944
rect 145524 72904 145530 72916
rect 145926 72904 145932 72916
rect 145984 72904 145990 72956
rect 149974 72768 149980 72820
rect 150032 72808 150038 72820
rect 304994 72808 305000 72820
rect 150032 72780 305000 72808
rect 150032 72768 150038 72780
rect 304994 72768 305000 72780
rect 305052 72768 305058 72820
rect 149698 72700 149704 72752
rect 149756 72740 149762 72752
rect 307754 72740 307760 72752
rect 149756 72712 307760 72740
rect 149756 72700 149762 72712
rect 307754 72700 307760 72712
rect 307812 72700 307818 72752
rect 149790 72632 149796 72684
rect 149848 72672 149854 72684
rect 311894 72672 311900 72684
rect 149848 72644 311900 72672
rect 149848 72632 149854 72644
rect 311894 72632 311900 72644
rect 311952 72632 311958 72684
rect 151354 72564 151360 72616
rect 151412 72604 151418 72616
rect 332594 72604 332600 72616
rect 151412 72576 332600 72604
rect 151412 72564 151418 72576
rect 332594 72564 332600 72576
rect 332652 72564 332658 72616
rect 154482 72496 154488 72548
rect 154540 72536 154546 72548
rect 340874 72536 340880 72548
rect 154540 72508 340880 72536
rect 154540 72496 154546 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 96614 72428 96620 72480
rect 96672 72468 96678 72480
rect 133138 72468 133144 72480
rect 96672 72440 133144 72468
rect 96672 72428 96678 72440
rect 133138 72428 133144 72440
rect 133196 72428 133202 72480
rect 158622 72428 158628 72480
rect 158680 72468 158686 72480
rect 368474 72468 368480 72480
rect 158680 72440 368480 72468
rect 158680 72428 158686 72440
rect 368474 72428 368480 72440
rect 368532 72428 368538 72480
rect 124766 72360 124772 72412
rect 124824 72400 124830 72412
rect 125410 72400 125416 72412
rect 124824 72372 125416 72400
rect 124824 72360 124830 72372
rect 125410 72360 125416 72372
rect 125468 72360 125474 72412
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 17310 71720 17316 71732
rect 3476 71692 17316 71720
rect 3476 71680 3482 71692
rect 17310 71680 17316 71692
rect 17368 71680 17374 71732
rect 139118 71476 139124 71528
rect 139176 71516 139182 71528
rect 171134 71516 171140 71528
rect 139176 71488 171140 71516
rect 139176 71476 139182 71488
rect 171134 71476 171140 71488
rect 171192 71476 171198 71528
rect 155126 71408 155132 71460
rect 155184 71448 155190 71460
rect 382274 71448 382280 71460
rect 155184 71420 382280 71448
rect 155184 71408 155190 71420
rect 382274 71408 382280 71420
rect 382332 71408 382338 71460
rect 157978 71340 157984 71392
rect 158036 71380 158042 71392
rect 408494 71380 408500 71392
rect 158036 71352 408500 71380
rect 158036 71340 158042 71352
rect 408494 71340 408500 71352
rect 408552 71340 408558 71392
rect 163406 71272 163412 71324
rect 163464 71312 163470 71324
rect 490006 71312 490012 71324
rect 163464 71284 490012 71312
rect 163464 71272 163470 71284
rect 490006 71272 490012 71284
rect 490064 71272 490070 71324
rect 164970 71204 164976 71256
rect 165028 71244 165034 71256
rect 507854 71244 507860 71256
rect 165028 71216 507860 71244
rect 165028 71204 165034 71216
rect 507854 71204 507860 71216
rect 507912 71204 507918 71256
rect 166534 71136 166540 71188
rect 166592 71176 166598 71188
rect 523034 71176 523040 71188
rect 166592 71148 523040 71176
rect 166592 71136 166598 71148
rect 523034 71136 523040 71148
rect 523092 71136 523098 71188
rect 168006 71068 168012 71120
rect 168064 71108 168070 71120
rect 536834 71108 536840 71120
rect 168064 71080 536840 71108
rect 168064 71068 168070 71080
rect 536834 71068 536840 71080
rect 536892 71068 536898 71120
rect 167914 71000 167920 71052
rect 167972 71040 167978 71052
rect 539594 71040 539600 71052
rect 167972 71012 539600 71040
rect 167972 71000 167978 71012
rect 539594 71000 539600 71012
rect 539652 71000 539658 71052
rect 137278 70456 137284 70508
rect 137336 70456 137342 70508
rect 137296 70428 137324 70456
rect 138750 70428 138756 70440
rect 137296 70400 138756 70428
rect 138750 70388 138756 70400
rect 138808 70388 138814 70440
rect 166350 69708 166356 69760
rect 166408 69748 166414 69760
rect 518894 69748 518900 69760
rect 166408 69720 518900 69748
rect 166408 69708 166414 69720
rect 518894 69708 518900 69720
rect 518952 69708 518958 69760
rect 169478 69640 169484 69692
rect 169536 69680 169542 69692
rect 564526 69680 564532 69692
rect 169536 69652 564532 69680
rect 169536 69640 169542 69652
rect 564526 69640 564532 69652
rect 564584 69640 564590 69692
rect 140038 68416 140044 68468
rect 140096 68456 140102 68468
rect 184934 68456 184940 68468
rect 140096 68428 184940 68456
rect 140096 68416 140102 68428
rect 184934 68416 184940 68428
rect 184992 68416 184998 68468
rect 159266 68348 159272 68400
rect 159324 68388 159330 68400
rect 218698 68388 218704 68400
rect 159324 68360 218704 68388
rect 159324 68348 159330 68360
rect 218698 68348 218704 68360
rect 218756 68348 218762 68400
rect 156966 68280 156972 68332
rect 157024 68320 157030 68332
rect 320174 68320 320180 68332
rect 157024 68292 320180 68320
rect 157024 68280 157030 68292
rect 320174 68280 320180 68292
rect 320232 68280 320238 68332
rect 138566 67532 138572 67584
rect 138624 67572 138630 67584
rect 140038 67572 140044 67584
rect 138624 67544 140044 67572
rect 138624 67532 138630 67544
rect 140038 67532 140044 67544
rect 140096 67532 140102 67584
rect 139946 67056 139952 67108
rect 140004 67096 140010 67108
rect 189074 67096 189080 67108
rect 140004 67068 189080 67096
rect 140004 67056 140010 67068
rect 189074 67056 189080 67068
rect 189132 67056 189138 67108
rect 157886 66988 157892 67040
rect 157944 67028 157950 67040
rect 412634 67028 412640 67040
rect 157944 67000 412640 67028
rect 157944 66988 157950 67000
rect 412634 66988 412640 67000
rect 412692 66988 412698 67040
rect 167638 66920 167644 66972
rect 167696 66960 167702 66972
rect 543734 66960 543740 66972
rect 167696 66932 543740 66960
rect 167696 66920 167702 66932
rect 543734 66920 543740 66932
rect 543792 66920 543798 66972
rect 170214 66852 170220 66904
rect 170272 66892 170278 66904
rect 569954 66892 569960 66904
rect 170272 66864 569960 66892
rect 170272 66852 170278 66864
rect 569954 66852 569960 66864
rect 570012 66852 570018 66904
rect 155678 65628 155684 65680
rect 155736 65668 155742 65680
rect 367094 65668 367100 65680
rect 155736 65640 367100 65668
rect 155736 65628 155742 65640
rect 367094 65628 367100 65640
rect 367152 65628 367158 65680
rect 166258 65560 166264 65612
rect 166316 65600 166322 65612
rect 525794 65600 525800 65612
rect 166316 65572 525800 65600
rect 166316 65560 166322 65572
rect 525794 65560 525800 65572
rect 525852 65560 525858 65612
rect 170122 65492 170128 65544
rect 170180 65532 170186 65544
rect 572714 65532 572720 65544
rect 170180 65504 572720 65532
rect 170180 65492 170186 65504
rect 572714 65492 572720 65504
rect 572772 65492 572778 65544
rect 152458 64472 152464 64524
rect 152516 64512 152522 64524
rect 338114 64512 338120 64524
rect 152516 64484 338120 64512
rect 152516 64472 152522 64484
rect 338114 64472 338120 64484
rect 338172 64472 338178 64524
rect 152550 64404 152556 64456
rect 152608 64444 152614 64456
rect 339494 64444 339500 64456
rect 152608 64416 339500 64444
rect 152608 64404 152614 64416
rect 339494 64404 339500 64416
rect 339552 64404 339558 64456
rect 156690 64336 156696 64388
rect 156748 64376 156754 64388
rect 390554 64376 390560 64388
rect 156748 64348 390560 64376
rect 156748 64336 156754 64348
rect 390554 64336 390560 64348
rect 390612 64336 390618 64388
rect 162026 64268 162032 64320
rect 162084 64308 162090 64320
rect 463694 64308 463700 64320
rect 162084 64280 463700 64308
rect 162084 64268 162090 64280
rect 463694 64268 463700 64280
rect 463752 64268 463758 64320
rect 163406 64200 163412 64252
rect 163464 64240 163470 64252
rect 487154 64240 487160 64252
rect 163464 64212 487160 64240
rect 163464 64200 163470 64212
rect 487154 64200 487160 64212
rect 487212 64200 487218 64252
rect 170030 64132 170036 64184
rect 170088 64172 170094 64184
rect 568574 64172 568580 64184
rect 170088 64144 568580 64172
rect 170088 64132 170094 64144
rect 568574 64132 568580 64144
rect 568632 64132 568638 64184
rect 142798 62976 142804 63028
rect 142856 63016 142862 63028
rect 224954 63016 224960 63028
rect 142856 62988 224960 63016
rect 142856 62976 142862 62988
rect 224954 62976 224960 62988
rect 225012 62976 225018 63028
rect 152366 62908 152372 62960
rect 152424 62948 152430 62960
rect 340966 62948 340972 62960
rect 152424 62920 340972 62948
rect 152424 62908 152430 62920
rect 340966 62908 340972 62920
rect 341024 62908 341030 62960
rect 161934 62840 161940 62892
rect 161992 62880 161998 62892
rect 465074 62880 465080 62892
rect 161992 62852 465080 62880
rect 161992 62840 161998 62852
rect 465074 62840 465080 62852
rect 465132 62840 465138 62892
rect 170490 62772 170496 62824
rect 170548 62812 170554 62824
rect 514754 62812 514760 62824
rect 170548 62784 514760 62812
rect 170548 62772 170554 62784
rect 514754 62772 514760 62784
rect 514812 62772 514818 62824
rect 149606 61412 149612 61464
rect 149664 61452 149670 61464
rect 303614 61452 303620 61464
rect 149664 61424 303620 61452
rect 149664 61412 149670 61424
rect 303614 61412 303620 61424
rect 303672 61412 303678 61464
rect 102226 61344 102232 61396
rect 102284 61384 102290 61396
rect 125318 61384 125324 61396
rect 102284 61356 125324 61384
rect 102284 61344 102290 61356
rect 125318 61344 125324 61356
rect 125376 61344 125382 61396
rect 138474 61344 138480 61396
rect 138532 61384 138538 61396
rect 152458 61384 152464 61396
rect 138532 61356 152464 61384
rect 138532 61344 138538 61356
rect 152458 61344 152464 61356
rect 152516 61344 152522 61396
rect 157794 61344 157800 61396
rect 157852 61384 157858 61396
rect 415394 61384 415400 61396
rect 157852 61356 415400 61384
rect 157852 61344 157858 61356
rect 415394 61344 415400 61356
rect 415452 61344 415458 61396
rect 182910 60664 182916 60716
rect 182968 60704 182974 60716
rect 580166 60704 580172 60716
rect 182968 60676 580172 60704
rect 182968 60664 182974 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 120074 60188 120080 60240
rect 120132 60228 120138 60240
rect 123570 60228 123576 60240
rect 120132 60200 123576 60228
rect 120132 60188 120138 60200
rect 123570 60188 123576 60200
rect 123628 60188 123634 60240
rect 151078 60188 151084 60240
rect 151136 60228 151142 60240
rect 331214 60228 331220 60240
rect 151136 60200 331220 60228
rect 151136 60188 151142 60200
rect 331214 60188 331220 60200
rect 331272 60188 331278 60240
rect 153746 60120 153752 60172
rect 153804 60160 153810 60172
rect 362954 60160 362960 60172
rect 153804 60132 362960 60160
rect 153804 60120 153810 60132
rect 362954 60120 362960 60132
rect 363012 60120 363018 60172
rect 156598 60052 156604 60104
rect 156656 60092 156662 60104
rect 396074 60092 396080 60104
rect 156656 60064 396080 60092
rect 156656 60052 156662 60064
rect 396074 60052 396080 60064
rect 396132 60052 396138 60104
rect 159174 59984 159180 60036
rect 159232 60024 159238 60036
rect 427814 60024 427820 60036
rect 159232 59996 427820 60024
rect 159232 59984 159238 59996
rect 427814 59984 427820 59996
rect 427872 59984 427878 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 180886 59344 180892 59356
rect 3108 59316 180892 59344
rect 3108 59304 3114 59316
rect 180886 59304 180892 59316
rect 180944 59304 180950 59356
rect 158346 58692 158352 58744
rect 158404 58732 158410 58744
rect 374086 58732 374092 58744
rect 158404 58704 374092 58732
rect 158404 58692 158410 58704
rect 374086 58692 374092 58704
rect 374144 58692 374150 58744
rect 159082 58624 159088 58676
rect 159140 58664 159146 58676
rect 440234 58664 440240 58676
rect 159140 58636 440240 58664
rect 159140 58624 159146 58636
rect 440234 58624 440240 58636
rect 440292 58624 440298 58676
rect 150986 57264 150992 57316
rect 151044 57304 151050 57316
rect 325694 57304 325700 57316
rect 151044 57276 325700 57304
rect 151044 57264 151050 57276
rect 325694 57264 325700 57276
rect 325752 57264 325758 57316
rect 95234 57196 95240 57248
rect 95292 57236 95298 57248
rect 125226 57236 125232 57248
rect 95292 57208 125232 57236
rect 95292 57196 95298 57208
rect 125226 57196 125232 57208
rect 125284 57196 125290 57248
rect 157702 57196 157708 57248
rect 157760 57236 157766 57248
rect 415486 57236 415492 57248
rect 157760 57208 415492 57236
rect 157760 57196 157766 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 88334 55836 88340 55888
rect 88392 55876 88398 55888
rect 125042 55876 125048 55888
rect 88392 55848 125048 55876
rect 88392 55836 88398 55848
rect 125042 55836 125048 55848
rect 125100 55836 125106 55888
rect 13814 51688 13820 51740
rect 13872 51728 13878 51740
rect 125134 51728 125140 51740
rect 13872 51700 125140 51728
rect 13872 51688 13878 51700
rect 125134 51688 125140 51700
rect 125192 51688 125198 51740
rect 153654 50396 153660 50448
rect 153712 50436 153718 50448
rect 357434 50436 357440 50448
rect 153712 50408 357440 50436
rect 153712 50396 153718 50408
rect 357434 50396 357440 50408
rect 357492 50396 357498 50448
rect 171686 50328 171692 50380
rect 171744 50368 171750 50380
rect 425054 50368 425060 50380
rect 171744 50340 425060 50368
rect 171744 50328 171750 50340
rect 425054 50328 425060 50340
rect 425112 50328 425118 50380
rect 171778 49036 171784 49088
rect 171836 49076 171842 49088
rect 418154 49076 418160 49088
rect 171836 49048 418160 49076
rect 171836 49036 171842 49048
rect 418154 49036 418160 49048
rect 418212 49036 418218 49088
rect 163314 48968 163320 49020
rect 163372 49008 163378 49020
rect 485774 49008 485780 49020
rect 163372 48980 485780 49008
rect 163372 48968 163378 48980
rect 485774 48968 485780 48980
rect 485832 48968 485838 49020
rect 118234 46860 118240 46912
rect 118292 46900 118298 46912
rect 580166 46900 580172 46912
rect 118292 46872 580172 46900
rect 118292 46860 118298 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 174078 45540 174084 45552
rect 3476 45512 174084 45540
rect 3476 45500 3482 45512
rect 174078 45500 174084 45512
rect 174136 45500 174142 45552
rect 67634 44956 67640 45008
rect 67692 44996 67698 45008
rect 130194 44996 130200 45008
rect 67692 44968 130200 44996
rect 67692 44956 67698 44968
rect 130194 44956 130200 44968
rect 130252 44956 130258 45008
rect 30374 44888 30380 44940
rect 30432 44928 30438 44940
rect 127526 44928 127532 44940
rect 30432 44900 127532 44928
rect 30432 44888 30438 44900
rect 127526 44888 127532 44900
rect 127584 44888 127590 44940
rect 27614 44820 27620 44872
rect 27672 44860 27678 44872
rect 127618 44860 127624 44872
rect 27672 44832 127624 44860
rect 27672 44820 27678 44832
rect 127618 44820 127624 44832
rect 127676 44820 127682 44872
rect 45554 37884 45560 37936
rect 45612 37924 45618 37936
rect 116578 37924 116584 37936
rect 45612 37896 116584 37924
rect 45612 37884 45618 37896
rect 116578 37884 116584 37896
rect 116636 37884 116642 37936
rect 7558 36524 7564 36576
rect 7616 36564 7622 36576
rect 124214 36564 124220 36576
rect 7616 36536 124220 36564
rect 7616 36524 7622 36536
rect 124214 36524 124220 36536
rect 124272 36524 124278 36576
rect 148410 35368 148416 35420
rect 148468 35408 148474 35420
rect 291194 35408 291200 35420
rect 148468 35380 291200 35408
rect 148468 35368 148474 35380
rect 291194 35368 291200 35380
rect 291252 35368 291258 35420
rect 159726 35300 159732 35352
rect 159784 35340 159790 35352
rect 382366 35340 382372 35352
rect 159784 35312 382372 35340
rect 159784 35300 159790 35312
rect 382366 35300 382372 35312
rect 382424 35300 382430 35352
rect 162486 35232 162492 35284
rect 162544 35272 162550 35284
rect 390646 35272 390652 35284
rect 162544 35244 390652 35272
rect 162544 35232 162550 35244
rect 390646 35232 390652 35244
rect 390704 35232 390710 35284
rect 38654 35164 38660 35216
rect 38712 35204 38718 35216
rect 122190 35204 122196 35216
rect 38712 35176 122196 35204
rect 38712 35164 38718 35176
rect 122190 35164 122196 35176
rect 122248 35164 122254 35216
rect 160738 35164 160744 35216
rect 160796 35204 160802 35216
rect 447134 35204 447140 35216
rect 160796 35176 447140 35204
rect 160796 35164 160802 35176
rect 447134 35164 447140 35176
rect 447192 35164 447198 35216
rect 142706 33804 142712 33856
rect 142764 33844 142770 33856
rect 219434 33844 219440 33856
rect 142764 33816 219440 33844
rect 142764 33804 142770 33816
rect 219434 33804 219440 33816
rect 219492 33804 219498 33856
rect 144270 33736 144276 33788
rect 144328 33776 144334 33788
rect 234614 33776 234620 33788
rect 144328 33748 234620 33776
rect 144328 33736 144334 33748
rect 234614 33736 234620 33748
rect 234672 33736 234678 33788
rect 173342 33056 173348 33108
rect 173400 33096 173406 33108
rect 580166 33096 580172 33108
rect 173400 33068 580172 33096
rect 173400 33056 173406 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 141418 32852 141424 32904
rect 141476 32892 141482 32904
rect 198734 32892 198740 32904
rect 141476 32864 198740 32892
rect 141476 32852 141482 32864
rect 198734 32852 198740 32864
rect 198792 32852 198798 32904
rect 141510 32784 141516 32836
rect 141568 32824 141574 32836
rect 201494 32824 201500 32836
rect 141568 32796 201500 32824
rect 141568 32784 141574 32796
rect 201494 32784 201500 32796
rect 201552 32784 201558 32836
rect 148226 32716 148232 32768
rect 148284 32756 148290 32768
rect 285674 32756 285680 32768
rect 148284 32728 285680 32756
rect 148284 32716 148290 32728
rect 285674 32716 285680 32728
rect 285732 32716 285738 32768
rect 148318 32648 148324 32700
rect 148376 32688 148382 32700
rect 287054 32688 287060 32700
rect 148376 32660 287060 32688
rect 148376 32648 148382 32660
rect 287054 32648 287060 32660
rect 287112 32648 287118 32700
rect 150894 32580 150900 32632
rect 150952 32620 150958 32632
rect 321554 32620 321560 32632
rect 150952 32592 321560 32620
rect 150952 32580 150958 32592
rect 321554 32580 321560 32592
rect 321612 32580 321618 32632
rect 3418 32512 3424 32564
rect 3476 32552 3482 32564
rect 7650 32552 7656 32564
rect 3476 32524 7656 32552
rect 3476 32512 3482 32524
rect 7650 32512 7656 32524
rect 7708 32512 7714 32564
rect 152182 32512 152188 32564
rect 152240 32552 152246 32564
rect 346394 32552 346400 32564
rect 152240 32524 346400 32552
rect 152240 32512 152246 32524
rect 346394 32512 346400 32524
rect 346452 32512 346458 32564
rect 152274 32444 152280 32496
rect 152332 32484 152338 32496
rect 349154 32484 349160 32496
rect 152332 32456 349160 32484
rect 152332 32444 152338 32456
rect 349154 32444 349160 32456
rect 349212 32444 349218 32496
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 120810 32416 120816 32428
rect 31812 32388 120816 32416
rect 31812 32376 31818 32388
rect 120810 32376 120816 32388
rect 120868 32376 120874 32428
rect 161842 32376 161848 32428
rect 161900 32416 161906 32428
rect 466454 32416 466460 32428
rect 161900 32388 466460 32416
rect 161900 32376 161906 32388
rect 466454 32376 466460 32388
rect 466512 32376 466518 32428
rect 304258 31152 304264 31204
rect 304316 31192 304322 31204
rect 465166 31192 465172 31204
rect 304316 31164 465172 31192
rect 304316 31152 304322 31164
rect 465166 31152 465172 31164
rect 465224 31152 465230 31204
rect 166166 31084 166172 31136
rect 166224 31124 166230 31136
rect 524414 31124 524420 31136
rect 166224 31096 524420 31124
rect 166224 31084 166230 31096
rect 524414 31084 524420 31096
rect 524472 31084 524478 31136
rect 167546 31016 167552 31068
rect 167604 31056 167610 31068
rect 535454 31056 535460 31068
rect 167604 31028 535460 31056
rect 167604 31016 167610 31028
rect 535454 31016 535460 31028
rect 535512 31016 535518 31068
rect 142614 29928 142620 29980
rect 142672 29968 142678 29980
rect 215294 29968 215300 29980
rect 142672 29940 215300 29968
rect 142672 29928 142678 29940
rect 215294 29928 215300 29940
rect 215352 29928 215358 29980
rect 156506 29860 156512 29912
rect 156564 29900 156570 29912
rect 391934 29900 391940 29912
rect 156564 29872 391940 29900
rect 156564 29860 156570 29872
rect 391934 29860 391940 29872
rect 391992 29860 391998 29912
rect 157518 29792 157524 29844
rect 157576 29832 157582 29844
rect 409874 29832 409880 29844
rect 157576 29804 409880 29832
rect 157576 29792 157582 29804
rect 409874 29792 409880 29804
rect 409932 29792 409938 29844
rect 157610 29724 157616 29776
rect 157668 29764 157674 29776
rect 416774 29764 416780 29776
rect 157668 29736 416780 29764
rect 157668 29724 157674 29736
rect 416774 29724 416780 29736
rect 416832 29724 416838 29776
rect 158990 29656 158996 29708
rect 159048 29696 159054 29708
rect 434714 29696 434720 29708
rect 159048 29668 434720 29696
rect 159048 29656 159054 29668
rect 434714 29656 434720 29668
rect 434772 29656 434778 29708
rect 167454 29588 167460 29640
rect 167512 29628 167518 29640
rect 542354 29628 542360 29640
rect 167512 29600 542360 29628
rect 167512 29588 167518 29600
rect 542354 29588 542360 29600
rect 542412 29588 542418 29640
rect 141326 28568 141332 28620
rect 141384 28608 141390 28620
rect 201586 28608 201592 28620
rect 141384 28580 201592 28608
rect 141384 28568 141390 28580
rect 201586 28568 201592 28580
rect 201644 28568 201650 28620
rect 141234 28500 141240 28552
rect 141292 28540 141298 28552
rect 204254 28540 204260 28552
rect 141292 28512 204260 28540
rect 141292 28500 141298 28512
rect 204254 28500 204260 28512
rect 204312 28500 204318 28552
rect 141142 28432 141148 28484
rect 141200 28472 141206 28484
rect 208394 28472 208400 28484
rect 141200 28444 208400 28472
rect 141200 28432 141206 28444
rect 208394 28432 208400 28444
rect 208452 28432 208458 28484
rect 154114 28364 154120 28416
rect 154172 28404 154178 28416
rect 332686 28404 332692 28416
rect 154172 28376 332692 28404
rect 154172 28364 154178 28376
rect 332686 28364 332692 28376
rect 332744 28364 332750 28416
rect 155034 28296 155040 28348
rect 155092 28336 155098 28348
rect 378134 28336 378140 28348
rect 155092 28308 378140 28336
rect 155092 28296 155098 28308
rect 378134 28296 378140 28308
rect 378192 28296 378198 28348
rect 160646 28228 160652 28280
rect 160704 28268 160710 28280
rect 454034 28268 454040 28280
rect 160704 28240 454040 28268
rect 160704 28228 160710 28240
rect 454034 28228 454040 28240
rect 454092 28228 454098 28280
rect 139762 27276 139768 27328
rect 139820 27316 139826 27328
rect 179414 27316 179420 27328
rect 139820 27288 179420 27316
rect 139820 27276 139826 27288
rect 179414 27276 179420 27288
rect 179472 27276 179478 27328
rect 139854 27208 139860 27260
rect 139912 27248 139918 27260
rect 183554 27248 183560 27260
rect 139912 27220 183560 27248
rect 139912 27208 139918 27220
rect 183554 27208 183560 27220
rect 183612 27208 183618 27260
rect 139670 27140 139676 27192
rect 139728 27180 139734 27192
rect 186314 27180 186320 27192
rect 139728 27152 186320 27180
rect 139728 27140 139734 27152
rect 186314 27140 186320 27152
rect 186372 27140 186378 27192
rect 142522 27072 142528 27124
rect 142580 27112 142586 27124
rect 218054 27112 218060 27124
rect 142580 27084 218060 27112
rect 142580 27072 142586 27084
rect 218054 27072 218060 27084
rect 218112 27072 218118 27124
rect 172238 27004 172244 27056
rect 172296 27044 172302 27056
rect 411254 27044 411260 27056
rect 172296 27016 411260 27044
rect 172296 27004 172302 27016
rect 411254 27004 411260 27016
rect 411312 27004 411318 27056
rect 156414 26936 156420 26988
rect 156472 26976 156478 26988
rect 398834 26976 398840 26988
rect 156472 26948 398840 26976
rect 156472 26936 156478 26948
rect 398834 26936 398840 26948
rect 398892 26936 398898 26988
rect 168926 26868 168932 26920
rect 168984 26908 168990 26920
rect 560294 26908 560300 26920
rect 168984 26880 560300 26908
rect 168984 26868 168990 26880
rect 560294 26868 560300 26880
rect 560352 26868 560358 26920
rect 140314 25916 140320 25968
rect 140372 25956 140378 25968
rect 176746 25956 176752 25968
rect 140372 25928 176752 25956
rect 140372 25916 140378 25928
rect 176746 25916 176752 25928
rect 176804 25916 176810 25968
rect 148134 25848 148140 25900
rect 148192 25888 148198 25900
rect 289814 25888 289820 25900
rect 148192 25860 289820 25888
rect 148192 25848 148198 25860
rect 289814 25848 289820 25860
rect 289872 25848 289878 25900
rect 157426 25780 157432 25832
rect 157484 25820 157490 25832
rect 414014 25820 414020 25832
rect 157484 25792 414020 25820
rect 157484 25780 157490 25792
rect 414014 25780 414020 25792
rect 414072 25780 414078 25832
rect 168742 25712 168748 25764
rect 168800 25752 168806 25764
rect 556154 25752 556160 25764
rect 168800 25724 556160 25752
rect 168800 25712 168806 25724
rect 556154 25712 556160 25724
rect 556212 25712 556218 25764
rect 168834 25644 168840 25696
rect 168892 25684 168898 25696
rect 563054 25684 563060 25696
rect 168892 25656 563060 25684
rect 168892 25644 168898 25656
rect 563054 25644 563060 25656
rect 563112 25644 563118 25696
rect 169846 25576 169852 25628
rect 169904 25616 169910 25628
rect 571334 25616 571340 25628
rect 169904 25588 571340 25616
rect 169904 25576 169910 25588
rect 571334 25576 571340 25588
rect 571392 25576 571398 25628
rect 169938 25508 169944 25560
rect 169996 25548 170002 25560
rect 572806 25548 572812 25560
rect 169996 25520 572812 25548
rect 169996 25508 170002 25520
rect 572806 25508 572812 25520
rect 572864 25508 572870 25560
rect 148042 24488 148048 24540
rect 148100 24528 148106 24540
rect 292574 24528 292580 24540
rect 148100 24500 292580 24528
rect 148100 24488 148106 24500
rect 292574 24488 292580 24500
rect 292632 24488 292638 24540
rect 167086 24420 167092 24472
rect 167144 24460 167150 24472
rect 534074 24460 534080 24472
rect 167144 24432 534080 24460
rect 167144 24420 167150 24432
rect 534074 24420 534080 24432
rect 534132 24420 534138 24472
rect 167270 24352 167276 24404
rect 167328 24392 167334 24404
rect 538214 24392 538220 24404
rect 167328 24364 538220 24392
rect 167328 24352 167334 24364
rect 538214 24352 538220 24364
rect 538272 24352 538278 24404
rect 167362 24284 167368 24336
rect 167420 24324 167426 24336
rect 540974 24324 540980 24336
rect 167420 24296 540980 24324
rect 167420 24284 167426 24296
rect 540974 24284 540980 24296
rect 541032 24284 541038 24336
rect 167178 24216 167184 24268
rect 167236 24256 167242 24268
rect 545114 24256 545120 24268
rect 167236 24228 545120 24256
rect 167236 24216 167242 24228
rect 545114 24216 545120 24228
rect 545172 24216 545178 24268
rect 168650 24148 168656 24200
rect 168708 24188 168714 24200
rect 552014 24188 552020 24200
rect 168708 24160 552020 24188
rect 168708 24148 168714 24160
rect 552014 24148 552020 24160
rect 552072 24148 552078 24200
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 181070 24120 181076 24132
rect 3384 24092 181076 24120
rect 3384 24080 3390 24092
rect 181070 24080 181076 24092
rect 181128 24080 181134 24132
rect 182818 24080 182824 24132
rect 182876 24120 182882 24132
rect 579614 24120 579620 24132
rect 182876 24092 579620 24120
rect 182876 24080 182882 24092
rect 579614 24080 579620 24092
rect 579672 24080 579678 24132
rect 3418 23128 3424 23180
rect 3476 23168 3482 23180
rect 173986 23168 173992 23180
rect 3476 23140 173992 23168
rect 3476 23128 3482 23140
rect 173986 23128 173992 23140
rect 174044 23128 174050 23180
rect 172146 23060 172152 23112
rect 172204 23100 172210 23112
rect 397454 23100 397460 23112
rect 172204 23072 397460 23100
rect 172204 23060 172210 23072
rect 397454 23060 397460 23072
rect 397512 23060 397518 23112
rect 161750 22992 161756 23044
rect 161808 23032 161814 23044
rect 467834 23032 467840 23044
rect 161808 23004 467840 23032
rect 161808 22992 161814 23004
rect 467834 22992 467840 23004
rect 467892 22992 467898 23044
rect 166074 22924 166080 22976
rect 166132 22964 166138 22976
rect 516134 22964 516140 22976
rect 166132 22936 516140 22964
rect 166132 22924 166138 22936
rect 516134 22924 516140 22936
rect 516192 22924 516198 22976
rect 165982 22856 165988 22908
rect 166040 22896 166046 22908
rect 520274 22896 520280 22908
rect 166040 22868 520280 22896
rect 166040 22856 166046 22868
rect 520274 22856 520280 22868
rect 520332 22856 520338 22908
rect 165890 22788 165896 22840
rect 165948 22828 165954 22840
rect 527174 22828 527180 22840
rect 165948 22800 527180 22828
rect 165948 22788 165954 22800
rect 527174 22788 527180 22800
rect 527232 22788 527238 22840
rect 118326 22720 118332 22772
rect 118384 22760 118390 22772
rect 580258 22760 580264 22772
rect 118384 22732 580264 22760
rect 118384 22720 118390 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 152090 21632 152096 21684
rect 152148 21672 152154 21684
rect 343634 21672 343640 21684
rect 152148 21644 343640 21672
rect 152148 21632 152154 21644
rect 343634 21632 343640 21644
rect 343692 21632 343698 21684
rect 172054 21564 172060 21616
rect 172112 21604 172118 21616
rect 440326 21604 440332 21616
rect 172112 21576 440332 21604
rect 172112 21564 172118 21576
rect 440326 21564 440332 21576
rect 440384 21564 440390 21616
rect 158898 21496 158904 21548
rect 158956 21536 158962 21548
rect 436094 21536 436100 21548
rect 158956 21508 436100 21536
rect 158956 21496 158962 21508
rect 436094 21496 436100 21508
rect 436152 21496 436158 21548
rect 163222 21428 163228 21480
rect 163280 21468 163286 21480
rect 484394 21468 484400 21480
rect 163280 21440 484400 21468
rect 163280 21428 163286 21440
rect 484394 21428 484400 21440
rect 484452 21428 484458 21480
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 126146 21400 126152 21412
rect 11112 21372 126152 21400
rect 11112 21360 11118 21372
rect 126146 21360 126152 21372
rect 126204 21360 126210 21412
rect 163130 21360 163136 21412
rect 163188 21400 163194 21412
rect 491294 21400 491300 21412
rect 163188 21372 491300 21400
rect 163188 21360 163194 21372
rect 491294 21360 491300 21372
rect 491352 21360 491358 21412
rect 145466 20612 145472 20664
rect 145524 20652 145530 20664
rect 262214 20652 262220 20664
rect 145524 20624 262220 20652
rect 145524 20612 145530 20624
rect 262214 20612 262220 20624
rect 262272 20612 262278 20664
rect 150802 20544 150808 20596
rect 150860 20584 150866 20596
rect 329834 20584 329840 20596
rect 150860 20556 329840 20584
rect 150860 20544 150866 20556
rect 329834 20544 329840 20556
rect 329892 20544 329898 20596
rect 145650 20476 145656 20528
rect 145708 20516 145714 20528
rect 255314 20516 255320 20528
rect 145708 20488 255320 20516
rect 145708 20476 145714 20488
rect 255314 20476 255320 20488
rect 255372 20476 255378 20528
rect 255958 20476 255964 20528
rect 256016 20516 256022 20528
rect 456886 20516 456892 20528
rect 256016 20488 456892 20516
rect 256016 20476 256022 20488
rect 456886 20476 456892 20488
rect 456944 20476 456950 20528
rect 242158 20408 242164 20460
rect 242216 20448 242222 20460
rect 449894 20448 449900 20460
rect 242216 20420 449900 20448
rect 242216 20408 242222 20420
rect 449894 20408 449900 20420
rect 449952 20408 449958 20460
rect 160278 20340 160284 20392
rect 160336 20380 160342 20392
rect 445754 20380 445760 20392
rect 160336 20352 445760 20380
rect 160336 20340 160342 20352
rect 445754 20340 445760 20352
rect 445812 20340 445818 20392
rect 160462 20272 160468 20324
rect 160520 20312 160526 20324
rect 448514 20312 448520 20324
rect 160520 20284 448520 20312
rect 160520 20272 160526 20284
rect 448514 20272 448520 20284
rect 448572 20272 448578 20324
rect 160186 20204 160192 20256
rect 160244 20244 160250 20256
rect 448606 20244 448612 20256
rect 160244 20216 448612 20244
rect 160244 20204 160250 20216
rect 448606 20204 448612 20216
rect 448664 20204 448670 20256
rect 160094 20136 160100 20188
rect 160152 20176 160158 20188
rect 451274 20176 451280 20188
rect 160152 20148 451280 20176
rect 160152 20136 160158 20148
rect 451274 20136 451280 20148
rect 451332 20136 451338 20188
rect 160554 20068 160560 20120
rect 160612 20108 160618 20120
rect 452654 20108 452660 20120
rect 160612 20080 452660 20108
rect 160612 20068 160618 20080
rect 452654 20068 452660 20080
rect 452712 20068 452718 20120
rect 160370 20000 160376 20052
rect 160428 20040 160434 20052
rect 455414 20040 455420 20052
rect 160428 20012 455420 20040
rect 160428 20000 160434 20012
rect 455414 20000 455420 20012
rect 455472 20000 455478 20052
rect 163038 19932 163044 19984
rect 163096 19972 163102 19984
rect 481726 19972 481732 19984
rect 163096 19944 481732 19972
rect 163096 19932 163102 19944
rect 481726 19932 481732 19944
rect 481784 19932 481790 19984
rect 145558 19864 145564 19916
rect 145616 19904 145622 19916
rect 259454 19904 259460 19916
rect 145616 19876 259460 19904
rect 145616 19864 145622 19876
rect 259454 19864 259460 19876
rect 259512 19864 259518 19916
rect 144178 18844 144184 18896
rect 144236 18884 144242 18896
rect 241514 18884 241520 18896
rect 144236 18856 241520 18884
rect 144236 18844 144242 18856
rect 241514 18844 241520 18856
rect 241572 18844 241578 18896
rect 171962 18776 171968 18828
rect 172020 18816 172026 18828
rect 404354 18816 404360 18828
rect 172020 18788 404360 18816
rect 172020 18776 172026 18788
rect 404354 18776 404360 18788
rect 404412 18776 404418 18828
rect 158806 18708 158812 18760
rect 158864 18748 158870 18760
rect 433334 18748 433340 18760
rect 158864 18720 433340 18748
rect 158864 18708 158870 18720
rect 433334 18708 433340 18720
rect 433392 18708 433398 18760
rect 63494 18640 63500 18692
rect 63552 18680 63558 18692
rect 126330 18680 126336 18692
rect 63552 18652 126336 18680
rect 63552 18640 63558 18652
rect 126330 18640 126336 18652
rect 126388 18640 126394 18692
rect 168466 18640 168472 18692
rect 168524 18680 168530 18692
rect 553394 18680 553400 18692
rect 168524 18652 553400 18680
rect 168524 18640 168530 18652
rect 553394 18640 553400 18652
rect 553452 18640 553458 18692
rect 42794 18572 42800 18624
rect 42852 18612 42858 18624
rect 128814 18612 128820 18624
rect 42852 18584 128820 18612
rect 42852 18572 42858 18584
rect 128814 18572 128820 18584
rect 128872 18572 128878 18624
rect 168558 18572 168564 18624
rect 168616 18612 168622 18624
rect 556246 18612 556252 18624
rect 168616 18584 556252 18612
rect 168616 18572 168622 18584
rect 556246 18572 556252 18584
rect 556304 18572 556310 18624
rect 142430 17824 142436 17876
rect 142488 17864 142494 17876
rect 216674 17864 216680 17876
rect 142488 17836 216680 17864
rect 142488 17824 142494 17836
rect 216674 17824 216680 17836
rect 216732 17824 216738 17876
rect 147122 17756 147128 17808
rect 147180 17796 147186 17808
rect 269114 17796 269120 17808
rect 147180 17768 269120 17796
rect 147180 17756 147186 17768
rect 269114 17756 269120 17768
rect 269172 17756 269178 17808
rect 147030 17688 147036 17740
rect 147088 17728 147094 17740
rect 273254 17728 273260 17740
rect 147088 17700 273260 17728
rect 147088 17688 147094 17700
rect 273254 17688 273260 17700
rect 273312 17688 273318 17740
rect 146938 17620 146944 17672
rect 146996 17660 147002 17672
rect 276014 17660 276020 17672
rect 146996 17632 276020 17660
rect 146996 17620 147002 17632
rect 276014 17620 276020 17632
rect 276072 17620 276078 17672
rect 172422 17552 172428 17604
rect 172480 17592 172486 17604
rect 347774 17592 347780 17604
rect 172480 17564 347780 17592
rect 172480 17552 172486 17564
rect 347774 17552 347780 17564
rect 347832 17552 347838 17604
rect 157334 17484 157340 17536
rect 157392 17524 157398 17536
rect 419534 17524 419540 17536
rect 157392 17496 419540 17524
rect 157392 17484 157398 17496
rect 419534 17484 419540 17496
rect 419592 17484 419598 17536
rect 160002 17416 160008 17468
rect 160060 17456 160066 17468
rect 441614 17456 441620 17468
rect 160060 17428 441620 17456
rect 160060 17416 160066 17428
rect 441614 17416 441620 17428
rect 441672 17416 441678 17468
rect 162946 17348 162952 17400
rect 163004 17388 163010 17400
rect 492674 17388 492680 17400
rect 163004 17360 492680 17388
rect 163004 17348 163010 17360
rect 492674 17348 492680 17360
rect 492732 17348 492738 17400
rect 164786 17280 164792 17332
rect 164844 17320 164850 17332
rect 503714 17320 503720 17332
rect 164844 17292 503720 17320
rect 164844 17280 164850 17292
rect 503714 17280 503720 17292
rect 503772 17280 503778 17332
rect 165522 17212 165528 17264
rect 165580 17252 165586 17264
rect 514846 17252 514852 17264
rect 165580 17224 514852 17252
rect 165580 17212 165586 17224
rect 514846 17212 514852 17224
rect 514904 17212 514910 17264
rect 144086 16192 144092 16244
rect 144144 16232 144150 16244
rect 237650 16232 237656 16244
rect 144144 16204 237656 16232
rect 144144 16192 144150 16204
rect 237650 16192 237656 16204
rect 237708 16192 237714 16244
rect 151998 16124 152004 16176
rect 152056 16164 152062 16176
rect 342898 16164 342904 16176
rect 152056 16136 342904 16164
rect 152056 16124 152062 16136
rect 342898 16124 342904 16136
rect 342956 16124 342962 16176
rect 153562 16056 153568 16108
rect 153620 16096 153626 16108
rect 361114 16096 361120 16108
rect 153620 16068 361120 16096
rect 153620 16056 153626 16068
rect 361114 16056 361120 16068
rect 361172 16056 361178 16108
rect 156322 15988 156328 16040
rect 156380 16028 156386 16040
rect 395338 16028 395344 16040
rect 156380 16000 395344 16028
rect 156380 15988 156386 16000
rect 395338 15988 395344 16000
rect 395396 15988 395402 16040
rect 156230 15920 156236 15972
rect 156288 15960 156294 15972
rect 398926 15960 398932 15972
rect 156288 15932 398932 15960
rect 156288 15920 156294 15932
rect 398926 15920 398932 15932
rect 398984 15920 398990 15972
rect 156138 15852 156144 15904
rect 156196 15892 156202 15904
rect 402514 15892 402520 15904
rect 156196 15864 402520 15892
rect 156196 15852 156202 15864
rect 402514 15852 402520 15864
rect 402572 15852 402578 15904
rect 145282 15104 145288 15156
rect 145340 15144 145346 15156
rect 254210 15144 254216 15156
rect 145340 15116 254216 15144
rect 145340 15104 145346 15116
rect 254210 15104 254216 15116
rect 254268 15104 254274 15156
rect 145374 15036 145380 15088
rect 145432 15076 145438 15088
rect 258258 15076 258264 15088
rect 145432 15048 258264 15076
rect 145432 15036 145438 15048
rect 258258 15036 258264 15048
rect 258316 15036 258322 15088
rect 146846 14968 146852 15020
rect 146904 15008 146910 15020
rect 268378 15008 268384 15020
rect 146904 14980 268384 15008
rect 146904 14968 146910 14980
rect 268378 14968 268384 14980
rect 268436 14968 268442 15020
rect 146754 14900 146760 14952
rect 146812 14940 146818 14952
rect 272426 14940 272432 14952
rect 146812 14912 272432 14940
rect 146812 14900 146818 14912
rect 272426 14900 272432 14912
rect 272484 14900 272490 14952
rect 149514 14832 149520 14884
rect 149572 14872 149578 14884
rect 311434 14872 311440 14884
rect 149572 14844 311440 14872
rect 149572 14832 149578 14844
rect 311434 14832 311440 14844
rect 311492 14832 311498 14884
rect 154942 14764 154948 14816
rect 155000 14804 155006 14816
rect 379514 14804 379520 14816
rect 155000 14776 379520 14804
rect 155000 14764 155006 14776
rect 379514 14764 379520 14776
rect 379572 14764 379578 14816
rect 154758 14696 154764 14748
rect 154816 14736 154822 14748
rect 381170 14736 381176 14748
rect 154816 14708 381176 14736
rect 154816 14696 154822 14708
rect 381170 14696 381176 14708
rect 381228 14696 381234 14748
rect 154666 14628 154672 14680
rect 154724 14668 154730 14680
rect 384298 14668 384304 14680
rect 154724 14640 384304 14668
rect 154724 14628 154730 14640
rect 384298 14628 384304 14640
rect 384356 14628 384362 14680
rect 154850 14560 154856 14612
rect 154908 14600 154914 14612
rect 386690 14600 386696 14612
rect 154908 14572 386696 14600
rect 154908 14560 154914 14572
rect 386690 14560 386696 14572
rect 386748 14560 386754 14612
rect 164694 14492 164700 14544
rect 164752 14532 164758 14544
rect 500586 14532 500592 14544
rect 164752 14504 500592 14532
rect 164752 14492 164758 14504
rect 500586 14492 500592 14504
rect 500644 14492 500650 14544
rect 165798 14424 165804 14476
rect 165856 14464 165862 14476
rect 523770 14464 523776 14476
rect 165856 14436 523776 14464
rect 165856 14424 165862 14436
rect 523770 14424 523776 14436
rect 523828 14424 523834 14476
rect 145190 14356 145196 14408
rect 145248 14396 145254 14408
rect 251266 14396 251272 14408
rect 145248 14368 251272 14396
rect 145248 14356 145254 14368
rect 251266 14356 251272 14368
rect 251324 14356 251330 14408
rect 139578 14288 139584 14340
rect 139636 14328 139642 14340
rect 188522 14328 188528 14340
rect 139636 14300 188528 14328
rect 139636 14288 139642 14300
rect 188522 14288 188528 14300
rect 188580 14288 188586 14340
rect 151906 13404 151912 13456
rect 151964 13444 151970 13456
rect 349246 13444 349252 13456
rect 151964 13416 349252 13444
rect 151964 13404 151970 13416
rect 349246 13404 349252 13416
rect 349304 13404 349310 13456
rect 153286 13336 153292 13388
rect 153344 13376 153350 13388
rect 357526 13376 357532 13388
rect 153344 13348 357532 13376
rect 153344 13336 153350 13348
rect 357526 13336 357532 13348
rect 357584 13336 357590 13388
rect 153470 13268 153476 13320
rect 153528 13308 153534 13320
rect 359458 13308 359464 13320
rect 153528 13280 359464 13308
rect 153528 13268 153534 13280
rect 359458 13268 359464 13280
rect 359516 13268 359522 13320
rect 155586 13200 155592 13252
rect 155644 13240 155650 13252
rect 361850 13240 361856 13252
rect 155644 13212 361856 13240
rect 155644 13200 155650 13212
rect 361850 13200 361856 13212
rect 361908 13200 361914 13252
rect 153378 13132 153384 13184
rect 153436 13172 153442 13184
rect 365806 13172 365812 13184
rect 153436 13144 365812 13172
rect 153436 13132 153442 13144
rect 365806 13132 365812 13144
rect 365864 13132 365870 13184
rect 162854 13064 162860 13116
rect 162912 13104 162918 13116
rect 488810 13104 488816 13116
rect 162912 13076 488816 13104
rect 162912 13064 162918 13076
rect 488810 13064 488816 13076
rect 488868 13064 488874 13116
rect 143902 12384 143908 12436
rect 143960 12424 143966 12436
rect 236546 12424 236552 12436
rect 143960 12396 236552 12424
rect 143960 12384 143966 12396
rect 236546 12384 236552 12396
rect 236604 12384 236610 12436
rect 146662 12316 146668 12368
rect 146720 12356 146726 12368
rect 276106 12356 276112 12368
rect 146720 12328 276112 12356
rect 146720 12316 146726 12328
rect 276106 12316 276112 12328
rect 276164 12316 276170 12368
rect 150710 12248 150716 12300
rect 150768 12288 150774 12300
rect 327994 12288 328000 12300
rect 150768 12260 328000 12288
rect 150768 12248 150774 12260
rect 327994 12248 328000 12260
rect 328052 12248 328058 12300
rect 150618 12180 150624 12232
rect 150676 12220 150682 12232
rect 328730 12220 328736 12232
rect 150676 12192 328736 12220
rect 150676 12180 150682 12192
rect 328730 12180 328736 12192
rect 328788 12180 328794 12232
rect 151814 12112 151820 12164
rect 151872 12152 151878 12164
rect 345290 12152 345296 12164
rect 151872 12124 345296 12152
rect 151872 12112 151878 12124
rect 345290 12112 345296 12124
rect 345348 12112 345354 12164
rect 156046 12044 156052 12096
rect 156104 12084 156110 12096
rect 400858 12084 400864 12096
rect 156104 12056 400864 12084
rect 156104 12044 156110 12056
rect 400858 12044 400864 12056
rect 400916 12044 400922 12096
rect 161658 11976 161664 12028
rect 161716 12016 161722 12028
rect 473446 12016 473452 12028
rect 161716 11988 473452 12016
rect 161716 11976 161722 11988
rect 473446 11976 473452 11988
rect 473504 11976 473510 12028
rect 164326 11908 164332 11960
rect 164384 11948 164390 11960
rect 498930 11948 498936 11960
rect 164384 11920 498936 11948
rect 164384 11908 164390 11920
rect 498930 11908 498936 11920
rect 498988 11908 498994 11960
rect 164418 11840 164424 11892
rect 164476 11880 164482 11892
rect 502978 11880 502984 11892
rect 164476 11852 502984 11880
rect 164476 11840 164482 11852
rect 502978 11840 502984 11852
rect 503036 11840 503042 11892
rect 117314 11772 117320 11824
rect 117372 11812 117378 11824
rect 134242 11812 134248 11824
rect 117372 11784 134248 11812
rect 117372 11772 117378 11784
rect 134242 11772 134248 11784
rect 134300 11772 134306 11824
rect 164510 11772 164516 11824
rect 164568 11812 164574 11824
rect 506474 11812 506480 11824
rect 164568 11784 506480 11812
rect 164568 11772 164574 11784
rect 506474 11772 506480 11784
rect 506532 11772 506538 11824
rect 106458 11704 106464 11756
rect 106516 11744 106522 11756
rect 133046 11744 133052 11756
rect 106516 11716 133052 11744
rect 106516 11704 106522 11716
rect 133046 11704 133052 11716
rect 133104 11704 133110 11756
rect 164602 11704 164608 11756
rect 164660 11744 164666 11756
rect 509602 11744 509608 11756
rect 164660 11716 509608 11744
rect 164660 11704 164666 11716
rect 509602 11704 509608 11716
rect 509660 11704 509666 11756
rect 143994 11636 144000 11688
rect 144052 11676 144058 11688
rect 233418 11676 233424 11688
rect 144052 11648 233424 11676
rect 144052 11636 144058 11648
rect 233418 11636 233424 11648
rect 233476 11636 233482 11688
rect 162394 11568 162400 11620
rect 162452 11608 162458 11620
rect 240134 11608 240140 11620
rect 162452 11580 240140 11608
rect 162452 11568 162458 11580
rect 240134 11568 240140 11580
rect 240192 11568 240198 11620
rect 139486 11500 139492 11552
rect 139544 11540 139550 11552
rect 139544 11512 180794 11540
rect 139544 11500 139550 11512
rect 176654 11432 176660 11484
rect 176712 11472 176718 11484
rect 177850 11472 177856 11484
rect 176712 11444 177856 11472
rect 176712 11432 176718 11444
rect 177850 11432 177856 11444
rect 177908 11432 177914 11484
rect 180766 11404 180794 11512
rect 184934 11500 184940 11552
rect 184992 11540 184998 11552
rect 186130 11540 186136 11552
rect 184992 11512 186136 11540
rect 184992 11500 184998 11512
rect 186130 11500 186136 11512
rect 186188 11500 186194 11552
rect 201494 11500 201500 11552
rect 201552 11540 201558 11552
rect 202690 11540 202696 11552
rect 201552 11512 202696 11540
rect 201552 11500 201558 11512
rect 202690 11500 202696 11512
rect 202748 11500 202754 11552
rect 184934 11404 184940 11416
rect 180766 11376 184940 11404
rect 184934 11364 184940 11376
rect 184992 11364 184998 11416
rect 85666 10548 85672 10600
rect 85724 10588 85730 10600
rect 131666 10588 131672 10600
rect 85724 10560 131672 10588
rect 85724 10548 85730 10560
rect 131666 10548 131672 10560
rect 131724 10548 131730 10600
rect 81618 10480 81624 10532
rect 81676 10520 81682 10532
rect 131758 10520 131764 10532
rect 81676 10492 131764 10520
rect 81676 10480 81682 10492
rect 131758 10480 131764 10492
rect 131816 10480 131822 10532
rect 78122 10412 78128 10464
rect 78180 10452 78186 10464
rect 128354 10452 128360 10464
rect 78180 10424 128360 10452
rect 78180 10412 78186 10424
rect 128354 10412 128360 10424
rect 128412 10412 128418 10464
rect 150526 10412 150532 10464
rect 150584 10452 150590 10464
rect 324406 10452 324412 10464
rect 150584 10424 324412 10452
rect 150584 10412 150590 10424
rect 324406 10412 324412 10424
rect 324464 10412 324470 10464
rect 25314 10344 25320 10396
rect 25372 10384 25378 10396
rect 93118 10384 93124 10396
rect 25372 10356 93124 10384
rect 25372 10344 25378 10356
rect 93118 10344 93124 10356
rect 93176 10344 93182 10396
rect 99834 10344 99840 10396
rect 99892 10384 99898 10396
rect 132954 10384 132960 10396
rect 99892 10356 132960 10384
rect 99892 10344 99898 10356
rect 132954 10344 132960 10356
rect 133012 10344 133018 10396
rect 161566 10344 161572 10396
rect 161624 10384 161630 10396
rect 469858 10384 469864 10396
rect 161624 10356 469864 10384
rect 161624 10344 161630 10356
rect 469858 10344 469864 10356
rect 469916 10344 469922 10396
rect 35986 10276 35992 10328
rect 36044 10316 36050 10328
rect 127434 10316 127440 10328
rect 36044 10288 127440 10316
rect 36044 10276 36050 10288
rect 127434 10276 127440 10288
rect 127492 10276 127498 10328
rect 166994 10276 167000 10328
rect 167052 10316 167058 10328
rect 539686 10316 539692 10328
rect 167052 10288 539692 10316
rect 167052 10276 167058 10288
rect 539686 10276 539692 10288
rect 539744 10276 539750 10328
rect 146570 9528 146576 9580
rect 146628 9568 146634 9580
rect 278314 9568 278320 9580
rect 146628 9540 278320 9568
rect 146628 9528 146634 9540
rect 278314 9528 278320 9540
rect 278372 9528 278378 9580
rect 147858 9460 147864 9512
rect 147916 9500 147922 9512
rect 288986 9500 288992 9512
rect 147916 9472 288992 9500
rect 147916 9460 147922 9472
rect 288986 9460 288992 9472
rect 289044 9460 289050 9512
rect 147950 9392 147956 9444
rect 148008 9432 148014 9444
rect 292574 9432 292580 9444
rect 148008 9404 292580 9432
rect 148008 9392 148014 9404
rect 292574 9392 292580 9404
rect 292632 9392 292638 9444
rect 147766 9324 147772 9376
rect 147824 9364 147830 9376
rect 296070 9364 296076 9376
rect 147824 9336 296076 9364
rect 147824 9324 147830 9336
rect 296070 9324 296076 9336
rect 296128 9324 296134 9376
rect 60826 9256 60832 9308
rect 60884 9296 60890 9308
rect 128998 9296 129004 9308
rect 60884 9268 129004 9296
rect 60884 9256 60890 9268
rect 128998 9256 129004 9268
rect 129056 9256 129062 9308
rect 149146 9256 149152 9308
rect 149204 9296 149210 9308
rect 303154 9296 303160 9308
rect 149204 9268 303160 9296
rect 149204 9256 149210 9268
rect 303154 9256 303160 9268
rect 303212 9256 303218 9308
rect 59630 9188 59636 9240
rect 59688 9228 59694 9240
rect 130102 9228 130108 9240
rect 59688 9200 130108 9228
rect 59688 9188 59694 9200
rect 130102 9188 130108 9200
rect 130160 9188 130166 9240
rect 149422 9188 149428 9240
rect 149480 9228 149486 9240
rect 306742 9228 306748 9240
rect 149480 9200 306748 9228
rect 149480 9188 149486 9200
rect 306742 9188 306748 9200
rect 306800 9188 306806 9240
rect 52546 9120 52552 9172
rect 52604 9160 52610 9172
rect 128630 9160 128636 9172
rect 52604 9132 128636 9160
rect 52604 9120 52610 9132
rect 128630 9120 128636 9132
rect 128688 9120 128694 9172
rect 149330 9120 149336 9172
rect 149388 9160 149394 9172
rect 310238 9160 310244 9172
rect 149388 9132 310244 9160
rect 149388 9120 149394 9132
rect 310238 9120 310244 9132
rect 310296 9120 310302 9172
rect 53742 9052 53748 9104
rect 53800 9092 53806 9104
rect 128538 9092 128544 9104
rect 53800 9064 128544 9092
rect 53800 9052 53806 9064
rect 128538 9052 128544 9064
rect 128596 9052 128602 9104
rect 149238 9052 149244 9104
rect 149296 9092 149302 9104
rect 313826 9092 313832 9104
rect 149296 9064 313832 9092
rect 149296 9052 149302 9064
rect 313826 9052 313832 9064
rect 313884 9052 313890 9104
rect 45462 8984 45468 9036
rect 45520 9024 45526 9036
rect 128722 9024 128728 9036
rect 45520 8996 128728 9024
rect 45520 8984 45526 8996
rect 128722 8984 128728 8996
rect 128780 8984 128786 9036
rect 165430 8984 165436 9036
rect 165488 9024 165494 9036
rect 507670 9024 507676 9036
rect 165488 8996 507676 9024
rect 165488 8984 165494 8996
rect 507670 8984 507676 8996
rect 507728 8984 507734 9036
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 126054 8956 126060 8968
rect 10008 8928 126060 8956
rect 10008 8916 10014 8928
rect 126054 8916 126060 8928
rect 126112 8916 126118 8968
rect 165706 8916 165712 8968
rect 165764 8956 165770 8968
rect 521838 8956 521844 8968
rect 165764 8928 521844 8956
rect 165764 8916 165770 8928
rect 521838 8916 521844 8928
rect 521896 8916 521902 8968
rect 116394 7964 116400 8016
rect 116452 8004 116458 8016
rect 134150 8004 134156 8016
rect 116452 7976 134156 8004
rect 116452 7964 116458 7976
rect 134150 7964 134156 7976
rect 134208 7964 134214 8016
rect 105722 7896 105728 7948
rect 105780 7936 105786 7948
rect 132770 7936 132776 7948
rect 105780 7908 132776 7936
rect 105780 7896 105786 7908
rect 132770 7896 132776 7908
rect 132828 7896 132834 7948
rect 98638 7828 98644 7880
rect 98696 7868 98702 7880
rect 132862 7868 132868 7880
rect 98696 7840 132868 7868
rect 98696 7828 98702 7840
rect 132862 7828 132868 7840
rect 132920 7828 132926 7880
rect 142246 7828 142252 7880
rect 142304 7868 142310 7880
rect 222746 7868 222752 7880
rect 142304 7840 222752 7868
rect 142304 7828 142310 7840
rect 222746 7828 222752 7840
rect 222804 7828 222810 7880
rect 84470 7760 84476 7812
rect 84528 7800 84534 7812
rect 131574 7800 131580 7812
rect 84528 7772 131580 7800
rect 84528 7760 84534 7772
rect 131574 7760 131580 7772
rect 131632 7760 131638 7812
rect 149054 7760 149060 7812
rect 149112 7800 149118 7812
rect 307938 7800 307944 7812
rect 149112 7772 307944 7800
rect 149112 7760 149118 7772
rect 307938 7760 307944 7772
rect 307996 7760 308002 7812
rect 48958 7692 48964 7744
rect 49016 7732 49022 7744
rect 129182 7732 129188 7744
rect 49016 7704 129188 7732
rect 49016 7692 49022 7704
rect 129182 7692 129188 7704
rect 129240 7692 129246 7744
rect 150434 7692 150440 7744
rect 150492 7732 150498 7744
rect 323302 7732 323308 7744
rect 150492 7704 323308 7732
rect 150492 7692 150498 7704
rect 323302 7692 323308 7704
rect 323360 7692 323366 7744
rect 34790 7624 34796 7676
rect 34848 7664 34854 7676
rect 127342 7664 127348 7676
rect 34848 7636 127348 7664
rect 34848 7624 34854 7636
rect 127342 7624 127348 7636
rect 127400 7624 127406 7676
rect 155862 7624 155868 7676
rect 155920 7664 155926 7676
rect 385954 7664 385960 7676
rect 155920 7636 385960 7664
rect 155920 7624 155926 7636
rect 385954 7624 385960 7636
rect 386012 7624 386018 7676
rect 24210 7556 24216 7608
rect 24268 7596 24274 7608
rect 122098 7596 122104 7608
rect 24268 7568 122104 7596
rect 24268 7556 24274 7568
rect 122098 7556 122104 7568
rect 122156 7556 122162 7608
rect 158714 7556 158720 7608
rect 158772 7596 158778 7608
rect 429654 7596 429660 7608
rect 158772 7568 429660 7596
rect 158772 7556 158778 7568
rect 429654 7556 429660 7568
rect 429712 7556 429718 7608
rect 139394 6808 139400 6860
rect 139452 6848 139458 6860
rect 181438 6848 181444 6860
rect 139452 6820 181444 6848
rect 139452 6808 139458 6820
rect 181438 6808 181444 6820
rect 181496 6808 181502 6860
rect 143810 6740 143816 6792
rect 143868 6780 143874 6792
rect 239306 6780 239312 6792
rect 143868 6752 239312 6780
rect 143868 6740 143874 6752
rect 239306 6740 239312 6752
rect 239364 6740 239370 6792
rect 143718 6672 143724 6724
rect 143776 6712 143782 6724
rect 242986 6712 242992 6724
rect 143776 6684 242992 6712
rect 143776 6672 143782 6684
rect 242986 6672 242992 6684
rect 243044 6672 243050 6724
rect 104526 6604 104532 6656
rect 104584 6644 104590 6656
rect 132678 6644 132684 6656
rect 104584 6616 132684 6644
rect 104584 6604 104590 6616
rect 132678 6604 132684 6616
rect 132736 6604 132742 6656
rect 145098 6604 145104 6656
rect 145156 6644 145162 6656
rect 253474 6644 253480 6656
rect 145156 6616 253480 6644
rect 145156 6604 145162 6616
rect 253474 6604 253480 6616
rect 253532 6604 253538 6656
rect 80882 6536 80888 6588
rect 80940 6576 80946 6588
rect 131390 6576 131396 6588
rect 80940 6548 131396 6576
rect 80940 6536 80946 6548
rect 131390 6536 131396 6548
rect 131448 6536 131454 6588
rect 144914 6536 144920 6588
rect 144972 6576 144978 6588
rect 257062 6576 257068 6588
rect 144972 6548 257068 6576
rect 144972 6536 144978 6548
rect 257062 6536 257068 6548
rect 257120 6536 257126 6588
rect 77386 6468 77392 6520
rect 77444 6508 77450 6520
rect 131482 6508 131488 6520
rect 77444 6480 131488 6508
rect 77444 6468 77450 6480
rect 131482 6468 131488 6480
rect 131540 6468 131546 6520
rect 145006 6468 145012 6520
rect 145064 6508 145070 6520
rect 260650 6508 260656 6520
rect 145064 6480 260656 6508
rect 145064 6468 145070 6480
rect 260650 6468 260656 6480
rect 260708 6468 260714 6520
rect 66714 6400 66720 6452
rect 66772 6440 66778 6452
rect 130010 6440 130016 6452
rect 66772 6412 130016 6440
rect 66772 6400 66778 6412
rect 130010 6400 130016 6412
rect 130068 6400 130074 6452
rect 146386 6400 146392 6452
rect 146444 6440 146450 6452
rect 271230 6440 271236 6452
rect 146444 6412 271236 6440
rect 146444 6400 146450 6412
rect 271230 6400 271236 6412
rect 271288 6400 271294 6452
rect 44266 6332 44272 6384
rect 44324 6372 44330 6384
rect 128906 6372 128912 6384
rect 44324 6344 128912 6372
rect 44324 6332 44330 6344
rect 128906 6332 128912 6344
rect 128964 6332 128970 6384
rect 146478 6332 146484 6384
rect 146536 6372 146542 6384
rect 274818 6372 274824 6384
rect 146536 6344 274824 6372
rect 146536 6332 146542 6344
rect 274818 6332 274824 6344
rect 274876 6332 274882 6384
rect 33594 6264 33600 6316
rect 33652 6304 33658 6316
rect 127250 6304 127256 6316
rect 33652 6276 127256 6304
rect 33652 6264 33658 6276
rect 127250 6264 127256 6276
rect 127308 6264 127314 6316
rect 137002 6264 137008 6316
rect 137060 6304 137066 6316
rect 149514 6304 149520 6316
rect 137060 6276 149520 6304
rect 137060 6264 137066 6276
rect 149514 6264 149520 6276
rect 149572 6264 149578 6316
rect 155954 6264 155960 6316
rect 156012 6304 156018 6316
rect 394234 6304 394240 6316
rect 156012 6276 394240 6304
rect 156012 6264 156018 6276
rect 394234 6264 394240 6276
rect 394292 6264 394298 6316
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 124950 6236 124956 6248
rect 19484 6208 124956 6236
rect 19484 6196 19490 6208
rect 124950 6196 124956 6208
rect 125008 6196 125014 6248
rect 137094 6196 137100 6248
rect 137152 6236 137158 6248
rect 154206 6236 154212 6248
rect 137152 6208 154212 6236
rect 137152 6196 137158 6208
rect 154206 6196 154212 6208
rect 154264 6196 154270 6248
rect 161474 6196 161480 6248
rect 161532 6236 161538 6248
rect 471054 6236 471060 6248
rect 161532 6208 471060 6236
rect 161532 6196 161538 6208
rect 471054 6196 471060 6208
rect 471112 6196 471118 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 125962 6168 125968 6180
rect 18288 6140 125968 6168
rect 18288 6128 18294 6140
rect 125962 6128 125968 6140
rect 126020 6128 126026 6180
rect 137186 6128 137192 6180
rect 137244 6168 137250 6180
rect 157794 6168 157800 6180
rect 137244 6140 157800 6168
rect 137244 6128 137250 6140
rect 157794 6128 157800 6140
rect 157852 6128 157858 6180
rect 168374 6128 168380 6180
rect 168432 6168 168438 6180
rect 562042 6168 562048 6180
rect 168432 6140 562048 6168
rect 168432 6128 168438 6140
rect 562042 6128 562048 6140
rect 562100 6128 562106 6180
rect 108298 5312 108304 5364
rect 108356 5352 108362 5364
rect 113818 5352 113824 5364
rect 108356 5324 113824 5352
rect 108356 5312 108362 5324
rect 113818 5312 113824 5324
rect 113876 5312 113882 5364
rect 114002 5312 114008 5364
rect 114060 5352 114066 5364
rect 134058 5352 134064 5364
rect 114060 5324 134064 5352
rect 114060 5312 114066 5324
rect 134058 5312 134064 5324
rect 134116 5312 134122 5364
rect 101030 5244 101036 5296
rect 101088 5284 101094 5296
rect 133138 5284 133144 5296
rect 101088 5256 133144 5284
rect 101088 5244 101094 5256
rect 133138 5244 133144 5256
rect 133196 5244 133202 5296
rect 93946 5176 93952 5228
rect 94004 5216 94010 5228
rect 133322 5216 133328 5228
rect 94004 5188 133328 5216
rect 94004 5176 94010 5188
rect 133322 5176 133328 5188
rect 133380 5176 133386 5228
rect 138106 5176 138112 5228
rect 138164 5216 138170 5228
rect 166074 5216 166080 5228
rect 138164 5188 166080 5216
rect 138164 5176 138170 5188
rect 166074 5176 166080 5188
rect 166132 5176 166138 5228
rect 63218 5108 63224 5160
rect 63276 5148 63282 5160
rect 129918 5148 129924 5160
rect 63276 5120 129924 5148
rect 63276 5108 63282 5120
rect 129918 5108 129924 5120
rect 129976 5108 129982 5160
rect 141050 5108 141056 5160
rect 141108 5148 141114 5160
rect 206186 5148 206192 5160
rect 141108 5120 206192 5148
rect 141108 5108 141114 5120
rect 206186 5108 206192 5120
rect 206244 5108 206250 5160
rect 30098 5040 30104 5092
rect 30156 5080 30162 5092
rect 127158 5080 127164 5092
rect 30156 5052 127164 5080
rect 30156 5040 30162 5052
rect 127158 5040 127164 5052
rect 127216 5040 127222 5092
rect 147674 5040 147680 5092
rect 147732 5080 147738 5092
rect 294874 5080 294880 5092
rect 147732 5052 294880 5080
rect 147732 5040 147738 5052
rect 294874 5040 294880 5052
rect 294932 5040 294938 5092
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 108298 5012 108304 5024
rect 15988 4984 108304 5012
rect 15988 4972 15994 4984
rect 108298 4972 108304 4984
rect 108356 4972 108362 5024
rect 136910 4972 136916 5024
rect 136968 5012 136974 5024
rect 145926 5012 145932 5024
rect 136968 4984 145932 5012
rect 136968 4972 136974 4984
rect 145926 4972 145932 4984
rect 145984 4972 145990 5024
rect 154390 4972 154396 5024
rect 154448 5012 154454 5024
rect 364610 5012 364616 5024
rect 154448 4984 364616 5012
rect 154448 4972 154454 4984
rect 364610 4972 364616 4984
rect 364668 4972 364674 5024
rect 436830 4972 436836 5024
rect 436888 5012 436894 5024
rect 436888 4984 451274 5012
rect 436888 4972 436894 4984
rect 28902 4904 28908 4956
rect 28960 4944 28966 4956
rect 127066 4944 127072 4956
rect 28960 4916 127072 4944
rect 28960 4904 28966 4916
rect 127066 4904 127072 4916
rect 127124 4904 127130 4956
rect 138382 4904 138388 4956
rect 138440 4944 138446 4956
rect 167178 4944 167184 4956
rect 138440 4916 167184 4944
rect 138440 4904 138446 4916
rect 167178 4904 167184 4916
rect 167236 4904 167242 4956
rect 175918 4904 175924 4956
rect 175976 4944 175982 4956
rect 433242 4944 433248 4956
rect 175976 4916 433248 4944
rect 175976 4904 175982 4916
rect 433242 4904 433248 4916
rect 433300 4904 433306 4956
rect 451246 4944 451274 4984
rect 479334 4944 479340 4956
rect 451246 4916 479340 4944
rect 479334 4904 479340 4916
rect 479392 4904 479398 4956
rect 6454 4836 6460 4888
rect 6512 4876 6518 4888
rect 10318 4876 10324 4888
rect 6512 4848 10324 4876
rect 6512 4836 6518 4848
rect 10318 4836 10324 4848
rect 10376 4836 10382 4888
rect 13538 4836 13544 4888
rect 13596 4876 13602 4888
rect 125778 4876 125784 4888
rect 13596 4848 125784 4876
rect 13596 4836 13602 4848
rect 125778 4836 125784 4848
rect 125836 4836 125842 4888
rect 138290 4836 138296 4888
rect 138348 4876 138354 4888
rect 169570 4876 169576 4888
rect 138348 4848 169576 4876
rect 138348 4836 138354 4848
rect 169570 4836 169576 4848
rect 169628 4836 169634 4888
rect 170674 4836 170680 4888
rect 170732 4876 170738 4888
rect 480530 4876 480536 4888
rect 170732 4848 480536 4876
rect 170732 4836 170738 4848
rect 480530 4836 480536 4848
rect 480588 4836 480594 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 125870 4808 125876 4820
rect 8812 4780 125876 4808
rect 8812 4768 8818 4780
rect 125870 4768 125876 4780
rect 125928 4768 125934 4820
rect 138198 4768 138204 4820
rect 138256 4808 138262 4820
rect 162486 4808 162492 4820
rect 138256 4780 162492 4808
rect 138256 4768 138262 4780
rect 162486 4768 162492 4780
rect 162544 4768 162550 4820
rect 166626 4768 166632 4820
rect 166684 4808 166690 4820
rect 518342 4808 518348 4820
rect 166684 4780 518348 4808
rect 166684 4768 166690 4780
rect 518342 4768 518348 4780
rect 518400 4768 518406 4820
rect 147030 4196 147036 4208
rect 146864 4168 147036 4196
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 122834 4088 122840 4140
rect 122892 4128 122898 4140
rect 123478 4128 123484 4140
rect 122892 4100 123484 4128
rect 122892 4088 122898 4100
rect 123478 4088 123484 4100
rect 123536 4088 123542 4140
rect 138842 4088 138848 4140
rect 138900 4128 138906 4140
rect 143534 4128 143540 4140
rect 138900 4100 143540 4128
rect 138900 4088 138906 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
rect 143626 4088 143632 4140
rect 143684 4128 143690 4140
rect 146864 4128 146892 4168
rect 147030 4156 147036 4168
rect 147088 4156 147094 4208
rect 143684 4100 146892 4128
rect 143684 4088 143690 4100
rect 146938 4088 146944 4140
rect 146996 4128 147002 4140
rect 151814 4128 151820 4140
rect 146996 4100 151820 4128
rect 146996 4088 147002 4100
rect 151814 4088 151820 4100
rect 151872 4088 151878 4140
rect 161106 4088 161112 4140
rect 161164 4128 161170 4140
rect 182542 4128 182548 4140
rect 161164 4100 182548 4128
rect 161164 4088 161170 4100
rect 182542 4088 182548 4100
rect 182600 4088 182606 4140
rect 218698 4088 218704 4140
rect 218756 4128 218762 4140
rect 219342 4128 219348 4140
rect 218756 4100 219348 4128
rect 218756 4088 218762 4100
rect 219342 4088 219348 4100
rect 219400 4088 219406 4140
rect 123110 4020 123116 4072
rect 123168 4060 123174 4072
rect 131206 4060 131212 4072
rect 123168 4032 131212 4060
rect 123168 4020 123174 4032
rect 131206 4020 131212 4032
rect 131264 4020 131270 4072
rect 136818 4020 136824 4072
rect 136876 4060 136882 4072
rect 150618 4060 150624 4072
rect 136876 4032 150624 4060
rect 136876 4020 136882 4032
rect 150618 4020 150624 4032
rect 150676 4020 150682 4072
rect 152458 4020 152464 4072
rect 152516 4060 152522 4072
rect 163682 4060 163688 4072
rect 152516 4032 163688 4060
rect 152516 4020 152522 4032
rect 163682 4020 163688 4032
rect 163740 4020 163746 4072
rect 171870 4020 171876 4072
rect 171928 4060 171934 4072
rect 196802 4060 196808 4072
rect 171928 4032 196808 4060
rect 171928 4020 171934 4032
rect 196802 4020 196808 4032
rect 196860 4020 196866 4072
rect 131850 3992 131856 4004
rect 123128 3964 131856 3992
rect 87966 3884 87972 3936
rect 88024 3924 88030 3936
rect 122834 3924 122840 3936
rect 88024 3896 122840 3924
rect 88024 3884 88030 3896
rect 122834 3884 122840 3896
rect 122892 3884 122898 3936
rect 86862 3816 86868 3868
rect 86920 3856 86926 3868
rect 123128 3856 123156 3964
rect 131850 3952 131856 3964
rect 131908 3952 131914 4004
rect 140130 3952 140136 4004
rect 140188 3992 140194 4004
rect 164878 3992 164884 4004
rect 140188 3964 164884 3992
rect 140188 3952 140194 3964
rect 164878 3952 164884 3964
rect 164936 3952 164942 4004
rect 173158 3952 173164 4004
rect 173216 3992 173222 4004
rect 212166 3992 212172 4004
rect 173216 3964 212172 3992
rect 173216 3952 173222 3964
rect 212166 3952 212172 3964
rect 212224 3952 212230 4004
rect 124674 3884 124680 3936
rect 124732 3924 124738 3936
rect 134518 3924 134524 3936
rect 124732 3896 134524 3924
rect 124732 3884 124738 3896
rect 134518 3884 134524 3896
rect 134576 3884 134582 3936
rect 140774 3884 140780 3936
rect 140832 3924 140838 3936
rect 200298 3924 200304 3936
rect 140832 3896 200304 3924
rect 140832 3884 140838 3896
rect 200298 3884 200304 3896
rect 200356 3884 200362 3936
rect 131298 3856 131304 3868
rect 86920 3828 123156 3856
rect 123220 3828 131304 3856
rect 86920 3816 86926 3828
rect 83274 3748 83280 3800
rect 83332 3788 83338 3800
rect 123110 3788 123116 3800
rect 83332 3760 123116 3788
rect 83332 3748 83338 3760
rect 123110 3748 123116 3760
rect 123168 3748 123174 3800
rect 79686 3680 79692 3732
rect 79744 3720 79750 3732
rect 123220 3720 123248 3828
rect 131298 3816 131304 3828
rect 131356 3816 131362 3868
rect 138750 3816 138756 3868
rect 138808 3856 138814 3868
rect 138808 3828 140360 3856
rect 138808 3816 138814 3828
rect 140332 3788 140360 3828
rect 140866 3816 140872 3868
rect 140924 3856 140930 3868
rect 203886 3856 203892 3868
rect 140924 3828 203892 3856
rect 140924 3816 140930 3828
rect 203886 3816 203892 3828
rect 203944 3816 203950 3868
rect 146938 3788 146944 3800
rect 140332 3760 146944 3788
rect 146938 3748 146944 3760
rect 146996 3748 147002 3800
rect 147030 3748 147036 3800
rect 147088 3788 147094 3800
rect 232222 3788 232228 3800
rect 147088 3760 232228 3788
rect 147088 3748 147094 3760
rect 232222 3748 232228 3760
rect 232280 3748 232286 3800
rect 251174 3748 251180 3800
rect 251232 3788 251238 3800
rect 252370 3788 252376 3800
rect 251232 3760 252376 3788
rect 251232 3748 251238 3760
rect 252370 3748 252376 3760
rect 252428 3748 252434 3800
rect 79744 3692 123248 3720
rect 79744 3680 79750 3692
rect 123294 3680 123300 3732
rect 123352 3720 123358 3732
rect 130654 3720 130660 3732
rect 123352 3692 130660 3720
rect 123352 3680 123358 3692
rect 130654 3680 130660 3692
rect 130712 3680 130718 3732
rect 135162 3680 135168 3732
rect 135220 3720 135226 3732
rect 135220 3692 140268 3720
rect 135220 3680 135226 3692
rect 69106 3612 69112 3664
rect 69164 3652 69170 3664
rect 126238 3652 126244 3664
rect 69164 3624 126244 3652
rect 69164 3612 69170 3624
rect 126238 3612 126244 3624
rect 126296 3612 126302 3664
rect 127066 3612 127072 3664
rect 127124 3652 127130 3664
rect 130286 3652 130292 3664
rect 127124 3624 130292 3652
rect 127124 3612 127130 3624
rect 130286 3612 130292 3624
rect 130344 3612 130350 3664
rect 136542 3612 136548 3664
rect 136600 3652 136606 3664
rect 140240 3652 140268 3692
rect 146294 3680 146300 3732
rect 146352 3720 146358 3732
rect 267734 3720 267740 3732
rect 146352 3692 267740 3720
rect 146352 3680 146358 3692
rect 267734 3680 267740 3692
rect 267792 3680 267798 3732
rect 276014 3680 276020 3732
rect 276072 3720 276078 3732
rect 276750 3720 276756 3732
rect 276072 3692 276756 3720
rect 276072 3680 276078 3692
rect 276750 3680 276756 3692
rect 276808 3680 276814 3732
rect 284294 3680 284300 3732
rect 284352 3720 284358 3732
rect 285030 3720 285036 3732
rect 284352 3692 285036 3720
rect 284352 3680 284358 3692
rect 285030 3680 285036 3692
rect 285088 3680 285094 3732
rect 161290 3652 161296 3664
rect 136600 3624 140176 3652
rect 140240 3624 161296 3652
rect 136600 3612 136606 3624
rect 35894 3544 35900 3596
rect 35952 3584 35958 3596
rect 36814 3584 36820 3596
rect 35952 3556 36820 3584
rect 35952 3544 35958 3556
rect 36814 3544 36820 3556
rect 36872 3544 36878 3596
rect 65518 3544 65524 3596
rect 65576 3584 65582 3596
rect 123294 3584 123300 3596
rect 65576 3556 123300 3584
rect 65576 3544 65582 3556
rect 123294 3544 123300 3556
rect 123352 3544 123358 3596
rect 126422 3584 126428 3596
rect 123404 3556 126428 3584
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 123404 3516 123432 3556
rect 126422 3544 126428 3556
rect 126480 3544 126486 3596
rect 129366 3544 129372 3596
rect 129424 3584 129430 3596
rect 130470 3584 130476 3596
rect 129424 3556 130476 3584
rect 129424 3544 129430 3556
rect 130470 3544 130476 3556
rect 130528 3544 130534 3596
rect 135438 3544 135444 3596
rect 135496 3584 135502 3596
rect 140038 3584 140044 3596
rect 135496 3556 140044 3584
rect 135496 3544 135502 3556
rect 140038 3544 140044 3556
rect 140096 3544 140102 3596
rect 17092 3488 123432 3516
rect 17092 3476 17098 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124858 3516 124864 3528
rect 123536 3488 124864 3516
rect 123536 3476 123542 3488
rect 124858 3476 124864 3488
rect 124916 3476 124922 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128170 3516 128176 3528
rect 127032 3488 128176 3516
rect 127032 3476 127038 3488
rect 128170 3476 128176 3488
rect 128228 3476 128234 3528
rect 135714 3476 135720 3528
rect 135772 3516 135778 3528
rect 138842 3516 138848 3528
rect 135772 3488 138848 3516
rect 135772 3476 135778 3488
rect 138842 3476 138848 3488
rect 138900 3476 138906 3528
rect 140148 3516 140176 3624
rect 161290 3612 161296 3624
rect 161348 3612 161354 3664
rect 163774 3612 163780 3664
rect 163832 3652 163838 3664
rect 324314 3652 324320 3664
rect 163832 3624 324320 3652
rect 163832 3612 163838 3624
rect 324314 3612 324320 3624
rect 324372 3612 324378 3664
rect 140958 3544 140964 3596
rect 141016 3584 141022 3596
rect 207382 3584 207388 3596
rect 141016 3556 207388 3584
rect 141016 3544 141022 3556
rect 207382 3544 207388 3556
rect 207440 3544 207446 3596
rect 218054 3544 218060 3596
rect 218112 3584 218118 3596
rect 219250 3584 219256 3596
rect 218112 3556 219256 3584
rect 218112 3544 218118 3556
rect 219250 3544 219256 3556
rect 219308 3544 219314 3596
rect 219342 3544 219348 3596
rect 219400 3584 219406 3596
rect 437934 3584 437940 3596
rect 219400 3556 437940 3584
rect 219400 3544 219406 3556
rect 437934 3544 437940 3556
rect 437992 3544 437998 3596
rect 440234 3544 440240 3596
rect 440292 3584 440298 3596
rect 441522 3584 441528 3596
rect 440292 3556 441528 3584
rect 440292 3544 440298 3556
rect 441522 3544 441528 3556
rect 441580 3544 441586 3596
rect 448606 3544 448612 3596
rect 448664 3584 448670 3596
rect 449802 3584 449808 3596
rect 448664 3556 449808 3584
rect 448664 3544 448670 3556
rect 449802 3544 449808 3556
rect 449860 3544 449866 3596
rect 456886 3544 456892 3596
rect 456944 3584 456950 3596
rect 458082 3584 458088 3596
rect 456944 3556 458088 3584
rect 456944 3544 456950 3556
rect 458082 3544 458088 3556
rect 458140 3544 458146 3596
rect 473998 3544 474004 3596
rect 474056 3584 474062 3596
rect 474056 3556 480254 3584
rect 474056 3544 474062 3556
rect 144730 3516 144736 3528
rect 140148 3488 144736 3516
rect 144730 3476 144736 3488
rect 144788 3476 144794 3528
rect 170766 3516 170772 3528
rect 146956 3488 170772 3516
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 125686 3448 125692 3460
rect 12400 3420 125692 3448
rect 12400 3408 12406 3420
rect 125686 3408 125692 3420
rect 125744 3408 125750 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 135898 3448 135904 3460
rect 131816 3420 135904 3448
rect 131816 3408 131822 3420
rect 135898 3408 135904 3420
rect 135956 3408 135962 3460
rect 140130 3408 140136 3460
rect 140188 3448 140194 3460
rect 146956 3448 146984 3488
rect 170766 3476 170772 3488
rect 170824 3476 170830 3528
rect 173250 3476 173256 3528
rect 173308 3516 173314 3528
rect 175458 3516 175464 3528
rect 173308 3488 175464 3516
rect 173308 3476 173314 3488
rect 175458 3476 175464 3488
rect 175516 3476 175522 3528
rect 462774 3516 462780 3528
rect 175568 3488 462780 3516
rect 168374 3448 168380 3460
rect 140188 3420 146984 3448
rect 147140 3420 168380 3448
rect 140188 3408 140194 3420
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 142982 3340 142988 3392
rect 143040 3380 143046 3392
rect 147030 3380 147036 3392
rect 143040 3352 147036 3380
rect 143040 3340 143046 3352
rect 147030 3340 147036 3352
rect 147088 3340 147094 3392
rect 139026 3272 139032 3324
rect 139084 3312 139090 3324
rect 147140 3312 147168 3420
rect 168374 3408 168380 3420
rect 168432 3408 168438 3460
rect 172330 3408 172336 3460
rect 172388 3448 172394 3460
rect 175568 3448 175596 3488
rect 462774 3476 462780 3488
rect 462832 3476 462838 3528
rect 465074 3476 465080 3528
rect 465132 3516 465138 3528
rect 465902 3516 465908 3528
rect 465132 3488 465908 3516
rect 465132 3476 465138 3488
rect 465902 3476 465908 3488
rect 465960 3476 465966 3528
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474182 3516 474188 3528
rect 473412 3488 474188 3516
rect 473412 3476 473418 3488
rect 474182 3476 474188 3488
rect 474240 3476 474246 3528
rect 480226 3516 480254 3556
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 574796 3556 576854 3584
rect 574796 3544 574802 3556
rect 495894 3516 495900 3528
rect 480226 3488 495900 3516
rect 495894 3476 495900 3488
rect 495952 3476 495958 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 172388 3420 175596 3448
rect 172388 3408 172394 3420
rect 180334 3408 180340 3460
rect 180392 3448 180398 3460
rect 475746 3448 475752 3460
rect 180392 3420 475752 3448
rect 180392 3408 180398 3420
rect 475746 3408 475752 3420
rect 475804 3408 475810 3460
rect 481634 3408 481640 3460
rect 481692 3448 481698 3460
rect 482462 3448 482468 3460
rect 481692 3420 482468 3448
rect 481692 3408 481698 3420
rect 482462 3408 482468 3420
rect 482520 3408 482526 3460
rect 576826 3448 576854 3556
rect 580994 3448 581000 3460
rect 576826 3420 581000 3448
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 147214 3340 147220 3392
rect 147272 3380 147278 3392
rect 155402 3380 155408 3392
rect 147272 3352 155408 3380
rect 147272 3340 147278 3352
rect 155402 3340 155408 3352
rect 155460 3340 155466 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365806 3340 365812 3392
rect 365864 3380 365870 3392
rect 367002 3380 367008 3392
rect 365864 3352 367008 3380
rect 365864 3340 365870 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 416682 3380 416688 3392
rect 415544 3352 416688 3380
rect 415544 3340 415550 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 139084 3284 147168 3312
rect 139084 3272 139090 3284
rect 137738 3204 137744 3256
rect 137796 3244 137802 3256
rect 147122 3244 147128 3256
rect 137796 3216 147128 3244
rect 137796 3204 137802 3216
rect 147122 3204 147128 3216
rect 147180 3204 147186 3256
rect 135806 3136 135812 3188
rect 135864 3176 135870 3188
rect 141234 3176 141240 3188
rect 135864 3148 141240 3176
rect 135864 3136 135870 3148
rect 141234 3136 141240 3148
rect 141292 3136 141298 3188
rect 144454 3136 144460 3188
rect 144512 3176 144518 3188
rect 153010 3176 153016 3188
rect 144512 3148 153016 3176
rect 144512 3136 144518 3148
rect 153010 3136 153016 3148
rect 153068 3136 153074 3188
rect 132954 3068 132960 3120
rect 133012 3108 133018 3120
rect 135530 3108 135536 3120
rect 133012 3080 135536 3108
rect 133012 3068 133018 3080
rect 135530 3068 135536 3080
rect 135588 3068 135594 3120
rect 136726 3068 136732 3120
rect 136784 3108 136790 3120
rect 148318 3108 148324 3120
rect 136784 3080 148324 3108
rect 136784 3068 136790 3080
rect 148318 3068 148324 3080
rect 148376 3068 148382 3120
rect 124122 3000 124128 3052
rect 124180 3040 124186 3052
rect 125870 3040 125876 3052
rect 124180 3012 125876 3040
rect 124180 3000 124186 3012
rect 125870 3000 125876 3012
rect 125928 3000 125934 3052
rect 135622 3000 135628 3052
rect 135680 3040 135686 3052
rect 137646 3040 137652 3052
rect 135680 3012 137652 3040
rect 135680 3000 135686 3012
rect 137646 3000 137652 3012
rect 137704 3000 137710 3052
rect 152734 2932 152740 2984
rect 152792 2972 152798 2984
rect 156598 2972 156604 2984
rect 152792 2944 156604 2972
rect 152792 2932 152798 2944
rect 156598 2932 156604 2944
rect 156656 2932 156662 2984
rect 349154 1504 349160 1556
rect 349212 1544 349218 1556
rect 350442 1544 350448 1556
rect 349212 1516 350448 1544
rect 349212 1504 349218 1516
rect 350442 1504 350448 1516
rect 350500 1504 350506 1556
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 45284 700408 45336 700460
rect 170312 700408 170364 700460
rect 364984 700408 365036 700460
rect 397644 700408 397696 700460
rect 405004 700408 405056 700460
rect 413652 700408 413704 700460
rect 44640 700340 44692 700392
rect 235172 700340 235224 700392
rect 283840 700340 283892 700392
rect 293960 700340 294012 700392
rect 348792 700340 348844 700392
rect 396448 700340 396500 700392
rect 403624 700340 403676 700392
rect 478512 700340 478564 700392
rect 44732 700272 44784 700324
rect 300124 700272 300176 700324
rect 332508 700272 332560 700324
rect 397552 700272 397604 700324
rect 400864 700272 400916 700324
rect 543464 700272 543516 700324
rect 198740 699660 198792 699712
rect 202788 699660 202840 699712
rect 258724 699660 258776 699712
rect 267648 699660 267700 699712
rect 398104 696940 398156 696992
rect 580172 696940 580224 696992
rect 187976 694764 188028 694816
rect 198740 694764 198792 694816
rect 293960 693404 294012 693456
rect 305644 693404 305696 693456
rect 185584 691364 185636 691416
rect 187976 691364 188028 691416
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 399484 683136 399536 683188
rect 580172 683136 580224 683188
rect 253940 681776 253992 681828
rect 258724 681776 258776 681828
rect 305644 679600 305696 679652
rect 322204 679600 322256 679652
rect 239404 678240 239456 678292
rect 253940 678240 253992 678292
rect 147772 678036 147824 678088
rect 153200 678036 153252 678088
rect 147036 675520 147088 675572
rect 147772 675520 147824 675572
rect 236644 671168 236696 671220
rect 239404 671168 239456 671220
rect 3516 670692 3568 670744
rect 18604 670692 18656 670744
rect 145564 667836 145616 667888
rect 147036 667836 147088 667888
rect 231308 662396 231360 662448
rect 236644 662396 236696 662448
rect 224224 659744 224276 659796
rect 231308 659744 231360 659796
rect 142804 657976 142856 658028
rect 145564 657976 145616 658028
rect 177856 653352 177908 653404
rect 185584 653352 185636 653404
rect 138388 652672 138440 652724
rect 142804 652740 142856 652792
rect 174820 646688 174872 646740
rect 177856 646688 177908 646740
rect 135904 644376 135956 644428
rect 138388 644444 138440 644496
rect 396724 643084 396776 643136
rect 580172 643084 580224 643136
rect 214564 638868 214616 638920
rect 218060 638868 218112 638920
rect 152464 638188 152516 638240
rect 174820 638188 174872 638240
rect 3516 632068 3568 632120
rect 7564 632068 7616 632120
rect 210424 632068 210476 632120
rect 214564 632068 214616 632120
rect 133144 630640 133196 630692
rect 135904 630640 135956 630692
rect 417424 630640 417476 630692
rect 579988 630640 580040 630692
rect 129740 623772 129792 623824
rect 133144 623772 133196 623824
rect 214564 623024 214616 623076
rect 224224 623024 224276 623076
rect 322204 622412 322256 622464
rect 324964 622412 325016 622464
rect 129004 620984 129056 621036
rect 129740 620984 129792 621036
rect 196624 620236 196676 620288
rect 214564 620236 214616 620288
rect 3516 618264 3568 618316
rect 21364 618264 21416 618316
rect 207020 611872 207072 611924
rect 210424 611872 210476 611924
rect 130384 609220 130436 609272
rect 207020 609220 207072 609272
rect 189080 605072 189132 605124
rect 196624 605072 196676 605124
rect 181444 600448 181496 600500
rect 189080 600448 189132 600500
rect 127624 598816 127676 598868
rect 130384 598816 130436 598868
rect 149336 594804 149388 594856
rect 152464 594804 152516 594856
rect 146944 592016 146996 592068
rect 149336 592016 149388 592068
rect 159364 589908 159416 589960
rect 181444 589908 181496 589960
rect 124864 581612 124916 581664
rect 127624 581612 127676 581664
rect 2780 579912 2832 579964
rect 4896 579912 4948 579964
rect 414664 576852 414716 576904
rect 580172 576852 580224 576904
rect 324964 570596 325016 570648
rect 329104 570596 329156 570648
rect 3056 565836 3108 565888
rect 31024 565836 31076 565888
rect 141424 565088 141476 565140
rect 146944 565088 146996 565140
rect 138020 554752 138072 554804
rect 141424 554752 141476 554804
rect 135904 550536 135956 550588
rect 138020 550536 138072 550588
rect 155224 542512 155276 542564
rect 159364 542512 159416 542564
rect 127624 540880 127676 540932
rect 129004 540880 129056 540932
rect 329104 532652 329156 532704
rect 331220 532652 331272 532704
rect 126244 529864 126296 529916
rect 127624 529864 127676 529916
rect 331220 529184 331272 529236
rect 341524 529184 341576 529236
rect 3516 527824 3568 527876
rect 8944 527824 8996 527876
rect 413284 524424 413336 524476
rect 580080 524424 580132 524476
rect 124220 520208 124272 520260
rect 126244 520208 126296 520260
rect 122104 518916 122156 518968
rect 124864 518916 124916 518968
rect 341524 517896 341576 517948
rect 343640 517896 343692 517948
rect 3516 514768 3568 514820
rect 32404 514768 32456 514820
rect 123484 514768 123536 514820
rect 124220 514768 124272 514820
rect 343640 513272 343692 513324
rect 347044 513272 347096 513324
rect 118976 511844 119028 511896
rect 122104 511844 122156 511896
rect 116032 507832 116084 507884
rect 118976 507832 119028 507884
rect 102784 502936 102836 502988
rect 116032 502936 116084 502988
rect 100024 498176 100076 498228
rect 102784 498176 102836 498228
rect 152464 480292 152516 480344
rect 155224 480292 155276 480344
rect 347044 476008 347096 476060
rect 353300 476008 353352 476060
rect 3516 474716 3568 474768
rect 13084 474716 13136 474768
rect 353300 472404 353352 472456
rect 356060 472404 356112 472456
rect 522304 470568 522356 470620
rect 580080 470568 580132 470620
rect 142804 468460 142856 468512
rect 152464 468460 152516 468512
rect 356060 467712 356112 467764
rect 359004 467712 359056 467764
rect 97264 464720 97316 464772
rect 100024 464720 100076 464772
rect 359004 464312 359056 464364
rect 370504 464312 370556 464364
rect 3516 462340 3568 462392
rect 22744 462340 22796 462392
rect 370504 459484 370556 459536
rect 376300 459484 376352 459536
rect 88984 458804 89036 458856
rect 97264 458804 97316 458856
rect 376300 456356 376352 456408
rect 381544 456356 381596 456408
rect 120724 453296 120776 453348
rect 142804 453296 142856 453348
rect 381544 437384 381596 437436
rect 384304 437384 384356 437436
rect 125508 425688 125560 425740
rect 135904 425688 135956 425740
rect 113824 422900 113876 422952
rect 125508 422900 125560 422952
rect 3332 422288 3384 422340
rect 10324 422288 10376 422340
rect 122104 420180 122156 420232
rect 123484 420180 123536 420232
rect 86224 419500 86276 419552
rect 88984 419500 89036 419552
rect 409144 418140 409196 418192
rect 580080 418140 580132 418192
rect 384304 415352 384356 415404
rect 387708 415352 387760 415404
rect 387708 411884 387760 411936
rect 396540 411884 396592 411936
rect 83464 410116 83516 410168
rect 86224 410116 86276 410168
rect 3332 409844 3384 409896
rect 28264 409844 28316 409896
rect 396816 404336 396868 404388
rect 580080 404336 580132 404388
rect 119344 401616 119396 401668
rect 122104 401616 122156 401668
rect 116584 398828 116636 398880
rect 119344 398828 119396 398880
rect 69664 396720 69716 396772
rect 136640 396720 136692 396772
rect 68284 384956 68336 385008
rect 69664 384956 69716 385008
rect 102048 384276 102100 384328
rect 113824 384276 113876 384328
rect 398196 378156 398248 378208
rect 580080 378156 580132 378208
rect 98644 377748 98696 377800
rect 102048 377748 102100 377800
rect 3332 371220 3384 371272
rect 14464 371220 14516 371272
rect 77944 371220 77996 371272
rect 83464 371220 83516 371272
rect 114928 370744 114980 370796
rect 116584 370744 116636 370796
rect 112444 367752 112496 367804
rect 114928 367752 114980 367804
rect 418804 364352 418856 364404
rect 579804 364352 579856 364404
rect 117320 362924 117372 362976
rect 120724 362924 120776 362976
rect 65432 358776 65484 358828
rect 68284 358776 68336 358828
rect 64144 358096 64196 358148
rect 65432 358096 65484 358148
rect 92480 358028 92532 358080
rect 98644 358028 98696 358080
rect 113180 357008 113232 357060
rect 117320 357008 117372 357060
rect 79324 355308 79376 355360
rect 92480 355308 92532 355360
rect 111064 353268 111116 353320
rect 112444 353268 112496 353320
rect 396908 351908 396960 351960
rect 580080 351908 580132 351960
rect 45836 349800 45888 349852
rect 77944 349800 77996 349852
rect 106924 348712 106976 348764
rect 113180 348712 113232 348764
rect 109776 343612 109828 343664
rect 111064 343612 111116 343664
rect 108304 340008 108356 340060
rect 109776 340008 109828 340060
rect 104532 338240 104584 338292
rect 106924 338240 106976 338292
rect 100760 335316 100812 335368
rect 104532 335316 104584 335368
rect 76564 333208 76616 333260
rect 100760 333208 100812 333260
rect 76656 329536 76708 329588
rect 79324 329536 79376 329588
rect 72424 321376 72476 321428
rect 76564 321376 76616 321428
rect 62764 319404 62816 319456
rect 64144 319404 64196 319456
rect 73804 318996 73856 319048
rect 76656 318996 76708 319048
rect 3148 318792 3200 318844
rect 26884 318792 26936 318844
rect 58624 315256 58676 315308
rect 72424 315256 72476 315308
rect 407764 311856 407816 311908
rect 579988 311856 580040 311908
rect 62856 305600 62908 305652
rect 108304 305600 108356 305652
rect 61476 299412 61528 299464
rect 62764 299412 62816 299464
rect 54484 298732 54536 298784
rect 58624 298732 58676 298784
rect 397000 298120 397052 298172
rect 579988 298120 580040 298172
rect 68284 295332 68336 295384
rect 73804 295332 73856 295384
rect 61200 294040 61252 294092
rect 62856 294040 62908 294092
rect 60004 293972 60056 294024
rect 61476 293972 61528 294024
rect 3240 292544 3292 292596
rect 11704 292544 11756 292596
rect 59544 289688 59596 289740
rect 61200 289688 61252 289740
rect 65708 285676 65760 285728
rect 68284 285676 68336 285728
rect 45744 284316 45796 284368
rect 54484 284316 54536 284368
rect 57336 284316 57388 284368
rect 59544 284316 59596 284368
rect 57980 282888 58032 282940
rect 60004 282888 60056 282940
rect 53104 280780 53156 280832
rect 57336 280780 57388 280832
rect 53840 278740 53892 278792
rect 57888 278740 57940 278792
rect 61384 277380 61436 277432
rect 65708 277380 65760 277432
rect 51724 276020 51776 276072
rect 53104 276020 53156 276072
rect 504364 271872 504416 271924
rect 579988 271872 580040 271924
rect 47584 271124 47636 271176
rect 53840 271124 53892 271176
rect 3148 266364 3200 266416
rect 17224 266364 17276 266416
rect 45652 263576 45704 263628
rect 47584 263576 47636 263628
rect 45192 261468 45244 261520
rect 61384 261468 61436 261520
rect 406384 258068 406436 258120
rect 579988 258068 580040 258120
rect 3240 253920 3292 253972
rect 25504 253920 25556 253972
rect 48228 253172 48280 253224
rect 51724 253172 51776 253224
rect 45560 249432 45612 249484
rect 48228 249432 48280 249484
rect 397092 244264 397144 244316
rect 579988 244264 580040 244316
rect 45468 241340 45520 241392
rect 45836 241340 45888 241392
rect 44916 240864 44968 240916
rect 71780 240864 71832 240916
rect 45008 240796 45060 240848
rect 88340 240796 88392 240848
rect 45100 240728 45152 240780
rect 104900 240728 104952 240780
rect 3240 240116 3292 240168
rect 44824 240116 44876 240168
rect 45468 239708 45520 239760
rect 45928 239708 45980 239760
rect 45376 238756 45428 238808
rect 45744 238756 45796 238808
rect 45836 233112 45888 233164
rect 45652 232908 45704 232960
rect 73804 232908 73856 232960
rect 116400 232364 116452 232416
rect 394792 232228 394844 232280
rect 396540 232228 396592 232280
rect 393964 231820 394016 231872
rect 579804 231820 579856 231872
rect 45376 231072 45428 231124
rect 50988 231072 51040 231124
rect 118608 231072 118660 231124
rect 397644 231072 397696 231124
rect 45192 230460 45244 230512
rect 46940 230460 46992 230512
rect 391940 230460 391992 230512
rect 394792 230460 394844 230512
rect 174544 229848 174596 229900
rect 176660 229848 176712 229900
rect 235264 228488 235316 228540
rect 266544 228488 266596 228540
rect 166264 228420 166316 228472
rect 296720 228420 296772 228472
rect 300124 228420 300176 228472
rect 356520 228420 356572 228472
rect 50988 228352 51040 228404
rect 58624 228352 58676 228404
rect 180064 228352 180116 228404
rect 580172 228352 580224 228404
rect 3240 227740 3292 227792
rect 40684 227740 40736 227792
rect 116400 227740 116452 227792
rect 122104 227740 122156 227792
rect 233884 227740 233936 227792
rect 236552 227740 236604 227792
rect 46940 227468 46992 227520
rect 50344 227468 50396 227520
rect 180156 226992 180208 227044
rect 580724 226992 580776 227044
rect 45652 224204 45704 224256
rect 48964 224204 49016 224256
rect 73804 224204 73856 224256
rect 77944 224204 77996 224256
rect 389824 223524 389876 223576
rect 391940 223524 391992 223576
rect 58624 219852 58676 219904
rect 64880 219852 64932 219904
rect 387800 218084 387852 218136
rect 389824 218084 389876 218136
rect 48964 218016 49016 218068
rect 211804 218016 211856 218068
rect 580172 218016 580224 218068
rect 51724 217948 51776 218000
rect 50344 216044 50396 216096
rect 65524 216044 65576 216096
rect 40684 215908 40736 215960
rect 164240 215908 164292 215960
rect 64880 215296 64932 215348
rect 68284 215296 68336 215348
rect 77944 215228 77996 215280
rect 86224 215228 86276 215280
rect 122104 214548 122156 214600
rect 135904 214548 135956 214600
rect 378324 214548 378376 214600
rect 387800 214548 387852 214600
rect 3240 213936 3292 213988
rect 90364 213936 90416 213988
rect 374920 212440 374972 212492
rect 378324 212508 378376 212560
rect 370504 209788 370556 209840
rect 374920 209788 374972 209840
rect 68284 207612 68336 207664
rect 88248 207612 88300 207664
rect 118700 205640 118752 205692
rect 580172 205640 580224 205692
rect 88248 203532 88300 203584
rect 112444 203532 112496 203584
rect 154856 202104 154908 202156
rect 235264 202104 235316 202156
rect 153200 200744 153252 200796
rect 233884 200744 233936 200796
rect 148968 199384 149020 199436
rect 207020 199384 207072 199436
rect 86224 199180 86276 199232
rect 88800 199180 88852 199232
rect 112444 198908 112496 198960
rect 115204 198908 115256 198960
rect 158904 197956 158956 198008
rect 386420 197956 386472 198008
rect 151084 197412 151136 197464
rect 153200 197412 153252 197464
rect 152740 197344 152792 197396
rect 154856 197344 154908 197396
rect 367744 197344 367796 197396
rect 370504 197344 370556 197396
rect 154488 196732 154540 196784
rect 166264 196732 166316 196784
rect 147956 196664 148008 196716
rect 174544 196664 174596 196716
rect 156144 196596 156196 196648
rect 327080 196596 327132 196648
rect 135904 196256 135956 196308
rect 138480 196256 138532 196308
rect 56600 195916 56652 195968
rect 138112 195916 138164 195968
rect 157524 195916 157576 195968
rect 300124 195916 300176 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 51724 195644 51776 195696
rect 53472 195644 53524 195696
rect 115940 194556 115992 194608
rect 140780 194556 140832 194608
rect 88800 194488 88852 194540
rect 91744 194488 91796 194540
rect 180248 191836 180300 191888
rect 579804 191836 579856 191888
rect 140780 190952 140832 191004
rect 53472 190544 53524 190596
rect 55864 190544 55916 190596
rect 140780 190476 140832 190528
rect 144736 190476 144788 190528
rect 149612 190476 149664 190528
rect 140688 190408 140740 190460
rect 165436 190340 165488 190392
rect 140780 190204 140832 190256
rect 165436 189048 165488 189100
rect 3148 187688 3200 187740
rect 119344 187688 119396 187740
rect 144460 180956 144512 181008
rect 146024 180956 146076 181008
rect 91744 180820 91796 180872
rect 95884 180820 95936 180872
rect 121460 180072 121512 180124
rect 136364 180072 136416 180124
rect 135996 178848 136048 178900
rect 136548 178848 136600 178900
rect 122840 178644 122892 178696
rect 136456 178644 136508 178696
rect 211896 178032 211948 178084
rect 579988 178032 580040 178084
rect 124220 177284 124272 177336
rect 135996 177284 136048 177336
rect 65524 177216 65576 177268
rect 72424 177216 72476 177268
rect 366364 176672 366416 176724
rect 367744 176672 367796 176724
rect 126980 176060 127032 176112
rect 136272 176060 136324 176112
rect 125600 175924 125652 175976
rect 136180 175924 136232 175976
rect 141608 175924 141660 175976
rect 149336 175992 149388 176044
rect 144460 175516 144512 175568
rect 149980 175516 150032 175568
rect 162492 175924 162544 175976
rect 154396 175380 154448 175432
rect 128360 175176 128412 175228
rect 136364 175176 136416 175228
rect 142068 174768 142120 174820
rect 141700 174700 141752 174752
rect 144092 174700 144144 174752
rect 145472 174700 145524 174752
rect 152464 174632 152516 174684
rect 156512 174632 156564 174684
rect 161480 174496 161532 174548
rect 167000 174292 167052 174344
rect 133880 173884 133932 173936
rect 137376 173884 137428 173936
rect 149336 172932 149388 172984
rect 151452 172932 151504 172984
rect 158444 172932 158496 172984
rect 159640 172932 159692 172984
rect 162492 172932 162544 172984
rect 165528 172932 165580 172984
rect 131120 172524 131172 172576
rect 136640 172524 136692 172576
rect 138020 172116 138072 172168
rect 140780 172116 140832 172168
rect 135260 171640 135312 171692
rect 138664 171640 138716 171692
rect 132500 171096 132552 171148
rect 136732 171096 136784 171148
rect 55864 169736 55916 169788
rect 60740 169668 60792 169720
rect 142436 166268 142488 166320
rect 142620 166268 142672 166320
rect 146484 166268 146536 166320
rect 147588 166268 147640 166320
rect 118516 165588 118568 165640
rect 580172 165588 580224 165640
rect 60740 163276 60792 163328
rect 66260 163276 66312 163328
rect 3148 162868 3200 162920
rect 86224 162868 86276 162920
rect 72424 156612 72476 156664
rect 79324 156612 79376 156664
rect 66260 155864 66312 155916
rect 67640 155864 67692 155916
rect 67640 153144 67692 153196
rect 72424 153144 72476 153196
rect 345664 151784 345716 151836
rect 580172 151784 580224 151836
rect 79324 149676 79376 149728
rect 87604 149676 87656 149728
rect 3332 149064 3384 149116
rect 179420 149064 179472 149116
rect 158444 148384 158496 148436
rect 164976 148384 165028 148436
rect 3056 148316 3108 148368
rect 180800 148316 180852 148368
rect 25504 146888 25556 146940
rect 182180 146888 182232 146940
rect 95884 146208 95936 146260
rect 101404 146208 101456 146260
rect 146576 143488 146628 143540
rect 148048 143488 148100 143540
rect 155224 143488 155276 143540
rect 160100 143488 160152 143540
rect 165436 143488 165488 143540
rect 169944 143488 169996 143540
rect 137744 143420 137796 143472
rect 139584 143420 139636 143472
rect 146484 143420 146536 143472
rect 149612 143420 149664 143472
rect 152464 143420 152516 143472
rect 157432 143420 157484 143472
rect 164976 143420 165028 143472
rect 168380 143420 168432 143472
rect 153476 143352 153528 143404
rect 158996 143352 159048 143404
rect 150532 143080 150584 143132
rect 154580 143080 154632 143132
rect 163596 143080 163648 143132
rect 174636 143080 174688 143132
rect 144460 143012 144512 143064
rect 160560 143012 160612 143064
rect 163504 143012 163556 143064
rect 145472 142944 145524 142996
rect 163688 142944 163740 142996
rect 164516 143012 164568 143064
rect 176200 143012 176252 143064
rect 178040 142944 178092 142996
rect 142528 142876 142580 142928
rect 173072 142876 173124 142928
rect 118332 142808 118384 142860
rect 396816 142808 396868 142860
rect 142068 142196 142120 142248
rect 142436 142196 142488 142248
rect 140688 142128 140740 142180
rect 142252 142128 142304 142180
rect 149520 142128 149572 142180
rect 152740 142128 152792 142180
rect 72424 141788 72476 141840
rect 179512 141788 179564 141840
rect 117872 141720 117924 141772
rect 397092 141720 397144 141772
rect 119160 141652 119212 141704
rect 429200 141652 429252 141704
rect 119252 141584 119304 141636
rect 494060 141584 494112 141636
rect 119068 141516 119120 141568
rect 558920 141516 558972 141568
rect 118976 141448 119028 141500
rect 580264 141448 580316 141500
rect 118884 141380 118936 141432
rect 580356 141380 580408 141432
rect 116768 140972 116820 141024
rect 182916 140972 182968 141024
rect 117136 140904 117188 140956
rect 182364 140904 182416 140956
rect 116676 140836 116728 140888
rect 182640 140836 182692 140888
rect 116952 140768 117004 140820
rect 182456 140768 182508 140820
rect 160100 140292 160152 140344
rect 180432 140292 180484 140344
rect 118148 140224 118200 140276
rect 397000 140224 397052 140276
rect 117964 140156 118016 140208
rect 396908 140156 396960 140208
rect 118792 140088 118844 140140
rect 580632 140088 580684 140140
rect 117780 140020 117832 140072
rect 580908 140020 580960 140072
rect 179512 139816 179564 139868
rect 180984 139816 181036 139868
rect 120540 139748 120592 139800
rect 182272 139748 182324 139800
rect 120632 139680 120684 139732
rect 182824 139680 182876 139732
rect 117228 139612 117280 139664
rect 183008 139612 183060 139664
rect 116400 139544 116452 139596
rect 182732 139544 182784 139596
rect 116860 139476 116912 139528
rect 182548 139476 182600 139528
rect 3240 139408 3292 139460
rect 179512 139408 179564 139460
rect 361580 138048 361632 138100
rect 366364 138048 366416 138100
rect 189724 137980 189776 138032
rect 580172 137980 580224 138032
rect 101404 137232 101456 137284
rect 106924 137232 106976 137284
rect 3332 136620 3384 136672
rect 116584 136620 116636 136672
rect 3148 136552 3200 136604
rect 117228 136552 117280 136604
rect 118424 136552 118476 136604
rect 23480 136484 23532 136536
rect 118240 136484 118292 136536
rect 360844 135260 360896 135312
rect 361580 135260 361632 135312
rect 18604 135192 18656 135244
rect 118424 135192 118476 135244
rect 117872 134852 117924 134904
rect 118424 134852 118476 134904
rect 21364 133832 21416 133884
rect 117136 133832 117188 133884
rect 31024 132404 31076 132456
rect 116952 132404 117004 132456
rect 32404 132336 32456 132388
rect 116860 132336 116912 132388
rect 359464 131112 359516 131164
rect 360844 131112 360896 131164
rect 22744 131044 22796 131096
rect 116676 131044 116728 131096
rect 115204 130364 115256 130416
rect 120724 130364 120776 130416
rect 28264 129684 28316 129736
rect 116400 129684 116452 129736
rect 117320 129684 117372 129736
rect 4068 128256 4120 128308
rect 116768 128256 116820 128308
rect 117320 128256 117372 128308
rect 90364 126216 90416 126268
rect 117320 126216 117372 126268
rect 180340 125604 180392 125656
rect 580172 125604 580224 125656
rect 7656 123428 7708 123480
rect 117780 123428 117832 123480
rect 17316 122068 17368 122120
rect 117688 122068 117740 122120
rect 106924 121456 106976 121508
rect 109684 121456 109736 121508
rect 86224 121388 86276 121440
rect 117320 121388 117372 121440
rect 180432 120776 180484 120828
rect 182180 120776 182232 120828
rect 6184 120096 6236 120148
rect 117412 120096 117464 120148
rect 17224 118600 17276 118652
rect 117320 118600 117372 118652
rect 87604 118532 87656 118584
rect 92480 118532 92532 118584
rect 14464 117240 14516 117292
rect 117412 117240 117464 117292
rect 26884 117172 26936 117224
rect 117320 117172 117372 117224
rect 10324 115880 10376 115932
rect 117320 115880 117372 115932
rect 92480 114520 92532 114572
rect 95884 114520 95936 114572
rect 13084 114452 13136 114504
rect 117320 114452 117372 114504
rect 8944 113092 8996 113144
rect 117320 113092 117372 113144
rect 180432 111800 180484 111852
rect 580172 111800 580224 111852
rect 4896 111732 4948 111784
rect 117320 111732 117372 111784
rect 7564 111664 7616 111716
rect 117412 111664 117464 111716
rect 3148 111460 3200 111512
rect 6184 111460 6236 111512
rect 357440 110440 357492 110492
rect 359464 110440 359516 110492
rect 4804 110372 4856 110424
rect 117320 110372 117372 110424
rect 182824 109692 182876 109744
rect 211804 109692 211856 109744
rect 40040 108944 40092 108996
rect 117320 108944 117372 108996
rect 45100 107584 45152 107636
rect 117320 107584 117372 107636
rect 183284 107584 183336 107636
rect 357440 107584 357492 107636
rect 45284 106224 45336 106276
rect 117320 106224 117372 106276
rect 183284 106224 183336 106276
rect 396448 106224 396500 106276
rect 44640 106156 44692 106208
rect 117412 106156 117464 106208
rect 44732 104796 44784 104848
rect 117320 104796 117372 104848
rect 183284 104796 183336 104848
rect 405004 104796 405056 104848
rect 95884 104728 95936 104780
rect 99564 104728 99616 104780
rect 183284 103436 183336 103488
rect 403624 103436 403676 103488
rect 183284 102076 183336 102128
rect 400864 102076 400916 102128
rect 109684 101396 109736 101448
rect 119436 101396 119488 101448
rect 183192 100648 183244 100700
rect 399484 100648 399536 100700
rect 238024 99356 238076 99408
rect 580172 99356 580224 99408
rect 183192 99288 183244 99340
rect 417424 99288 417476 99340
rect 99564 97928 99616 97980
rect 102784 97928 102836 97980
rect 183192 97928 183244 97980
rect 414664 97928 414716 97980
rect 183192 96568 183244 96620
rect 413284 96568 413336 96620
rect 183468 95140 183520 95192
rect 522304 95140 522356 95192
rect 183468 93780 183520 93832
rect 409144 93780 409196 93832
rect 183468 92420 183520 92472
rect 418804 92420 418856 92472
rect 102784 90992 102836 91044
rect 105636 90992 105688 91044
rect 183468 90992 183520 91044
rect 407764 90992 407816 91044
rect 182272 89632 182324 89684
rect 406384 89632 406436 89684
rect 182732 87592 182784 87644
rect 211896 87592 211948 87644
rect 105636 86912 105688 86964
rect 108120 86912 108172 86964
rect 179972 85552 180024 85604
rect 580172 85552 580224 85604
rect 182732 85484 182784 85536
rect 189724 85484 189776 85536
rect 3148 84192 3200 84244
rect 120632 84192 120684 84244
rect 182732 84124 182784 84176
rect 238024 84124 238076 84176
rect 178960 81200 179012 81252
rect 180340 81200 180392 81252
rect 108120 80724 108172 80776
rect 120080 80724 120132 80776
rect 178960 80724 179012 80776
rect 118516 80588 118568 80640
rect 118608 80520 118660 80572
rect 174452 80520 174504 80572
rect 178592 80656 178644 80708
rect 179972 80656 180024 80708
rect 174452 80384 174504 80436
rect 175280 80384 175332 80436
rect 345664 80724 345716 80776
rect 11704 79976 11756 80028
rect 3884 79840 3936 79892
rect 3700 79704 3752 79756
rect 3516 79568 3568 79620
rect 116584 79092 116636 79144
rect 123668 79840 123720 79892
rect 125738 79908 125790 79960
rect 126014 79908 126066 79960
rect 125508 79840 125560 79892
rect 125830 79840 125882 79892
rect 125048 79772 125100 79824
rect 125140 79636 125192 79688
rect 126198 79908 126250 79960
rect 126290 79908 126342 79960
rect 126382 79908 126434 79960
rect 126474 79908 126526 79960
rect 126658 79908 126710 79960
rect 126842 79908 126894 79960
rect 125876 79568 125928 79620
rect 126290 79772 126342 79824
rect 126336 79636 126388 79688
rect 125692 79432 125744 79484
rect 126704 79772 126756 79824
rect 127210 79840 127262 79892
rect 127026 79772 127078 79824
rect 126796 79704 126848 79756
rect 127486 79908 127538 79960
rect 127854 79908 127906 79960
rect 127946 79908 127998 79960
rect 128222 79908 128274 79960
rect 128406 79908 128458 79960
rect 128498 79908 128550 79960
rect 129050 79908 129102 79960
rect 129142 79908 129194 79960
rect 129510 79908 129562 79960
rect 129602 79908 129654 79960
rect 130154 79908 130206 79960
rect 130246 79908 130298 79960
rect 130706 79908 130758 79960
rect 130890 79908 130942 79960
rect 130982 79908 131034 79960
rect 131074 79908 131126 79960
rect 127394 79772 127446 79824
rect 127164 79704 127216 79756
rect 127256 79704 127308 79756
rect 127532 79704 127584 79756
rect 127808 79704 127860 79756
rect 127072 79636 127124 79688
rect 127348 79636 127400 79688
rect 128130 79840 128182 79892
rect 128176 79704 128228 79756
rect 128360 79704 128412 79756
rect 128590 79840 128642 79892
rect 128866 79840 128918 79892
rect 128774 79772 128826 79824
rect 128452 79636 128504 79688
rect 128544 79636 128596 79688
rect 128728 79636 128780 79688
rect 128958 79772 129010 79824
rect 128820 79568 128872 79620
rect 129326 79840 129378 79892
rect 129188 79772 129240 79824
rect 129096 79636 129148 79688
rect 129280 79636 129332 79688
rect 127624 79432 127676 79484
rect 128912 79500 128964 79552
rect 129004 79432 129056 79484
rect 129786 79840 129838 79892
rect 129970 79772 130022 79824
rect 130108 79772 130160 79824
rect 129740 79636 129792 79688
rect 130016 79636 130068 79688
rect 129556 79568 129608 79620
rect 130430 79840 130482 79892
rect 130614 79840 130666 79892
rect 129832 79500 129884 79552
rect 129924 79432 129976 79484
rect 130798 79840 130850 79892
rect 130660 79636 130712 79688
rect 130568 79568 130620 79620
rect 130292 79364 130344 79416
rect 130890 79772 130942 79824
rect 130936 79636 130988 79688
rect 131258 79908 131310 79960
rect 131442 79908 131494 79960
rect 131534 79908 131586 79960
rect 131626 79908 131678 79960
rect 131810 79908 131862 79960
rect 132270 79908 132322 79960
rect 132362 79908 132414 79960
rect 132454 79908 132506 79960
rect 132822 79908 132874 79960
rect 131304 79704 131356 79756
rect 131212 79636 131264 79688
rect 131580 79772 131632 79824
rect 131120 79568 131172 79620
rect 131488 79568 131540 79620
rect 132086 79840 132138 79892
rect 131994 79772 132046 79824
rect 132224 79704 132276 79756
rect 132638 79840 132690 79892
rect 132730 79840 132782 79892
rect 132592 79704 132644 79756
rect 132040 79636 132092 79688
rect 132132 79636 132184 79688
rect 132316 79636 132368 79688
rect 132684 79636 132736 79688
rect 133190 79908 133242 79960
rect 133650 79908 133702 79960
rect 133098 79840 133150 79892
rect 133466 79840 133518 79892
rect 133144 79704 133196 79756
rect 131948 79568 132000 79620
rect 133052 79568 133104 79620
rect 132684 79500 132736 79552
rect 133604 79636 133656 79688
rect 133512 79364 133564 79416
rect 134018 79908 134070 79960
rect 134570 79908 134622 79960
rect 134202 79840 134254 79892
rect 134386 79840 134438 79892
rect 133972 79772 134024 79824
rect 134110 79772 134162 79824
rect 134064 79568 134116 79620
rect 134248 79568 134300 79620
rect 134156 79500 134208 79552
rect 134524 79704 134576 79756
rect 134846 79908 134898 79960
rect 135214 79908 135266 79960
rect 135490 79908 135542 79960
rect 135582 79908 135634 79960
rect 135858 79908 135910 79960
rect 136226 79908 136278 79960
rect 136318 79908 136370 79960
rect 136410 79908 136462 79960
rect 136594 79908 136646 79960
rect 137054 79908 137106 79960
rect 135030 79840 135082 79892
rect 134616 79636 134668 79688
rect 134708 79636 134760 79688
rect 135306 79840 135358 79892
rect 135352 79704 135404 79756
rect 135444 79704 135496 79756
rect 135076 79568 135128 79620
rect 135260 79568 135312 79620
rect 135766 79772 135818 79824
rect 135720 79636 135772 79688
rect 136042 79840 136094 79892
rect 135904 79636 135956 79688
rect 135628 79500 135680 79552
rect 136686 79772 136738 79824
rect 136364 79704 136416 79756
rect 136180 79636 136232 79688
rect 136272 79636 136324 79688
rect 137606 79908 137658 79960
rect 137698 79908 137750 79960
rect 137974 79908 138026 79960
rect 137330 79840 137382 79892
rect 136824 79636 136876 79688
rect 136824 79500 136876 79552
rect 137284 79636 137336 79688
rect 137790 79840 137842 79892
rect 137652 79500 137704 79552
rect 137744 79500 137796 79552
rect 138250 79908 138302 79960
rect 138342 79908 138394 79960
rect 138526 79908 138578 79960
rect 138618 79908 138670 79960
rect 138710 79908 138762 79960
rect 138986 79908 139038 79960
rect 139170 79908 139222 79960
rect 138388 79636 138440 79688
rect 138480 79636 138532 79688
rect 138112 79568 138164 79620
rect 138296 79568 138348 79620
rect 138802 79840 138854 79892
rect 138894 79840 138946 79892
rect 138664 79704 138716 79756
rect 138756 79704 138808 79756
rect 139124 79772 139176 79824
rect 138940 79704 138992 79756
rect 139032 79704 139084 79756
rect 139032 79500 139084 79552
rect 139630 79908 139682 79960
rect 139722 79908 139774 79960
rect 139814 79908 139866 79960
rect 139906 79908 139958 79960
rect 139998 79908 140050 79960
rect 140182 79908 140234 79960
rect 140274 79908 140326 79960
rect 140366 79908 140418 79960
rect 140458 79908 140510 79960
rect 139538 79840 139590 79892
rect 139584 79704 139636 79756
rect 139676 79704 139728 79756
rect 139860 79704 139912 79756
rect 139768 79636 139820 79688
rect 140228 79772 140280 79824
rect 140826 79840 140878 79892
rect 140412 79772 140464 79824
rect 140136 79704 140188 79756
rect 140320 79636 140372 79688
rect 139584 79500 139636 79552
rect 141102 79772 141154 79824
rect 140872 79636 140924 79688
rect 141148 79636 141200 79688
rect 141470 79908 141522 79960
rect 141654 79908 141706 79960
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 141240 79568 141292 79620
rect 141056 79500 141108 79552
rect 138848 79432 138900 79484
rect 140964 79432 141016 79484
rect 141700 79772 141752 79824
rect 142022 79840 142074 79892
rect 141884 79704 141936 79756
rect 141792 79636 141844 79688
rect 142206 79908 142258 79960
rect 142298 79908 142350 79960
rect 143494 79908 143546 79960
rect 144874 79908 144926 79960
rect 144966 79908 145018 79960
rect 145058 79908 145110 79960
rect 145150 79908 145202 79960
rect 145242 79908 145294 79960
rect 142068 79704 142120 79756
rect 142666 79840 142718 79892
rect 142758 79840 142810 79892
rect 143218 79840 143270 79892
rect 143586 79840 143638 79892
rect 143770 79840 143822 79892
rect 144046 79840 144098 79892
rect 144322 79840 144374 79892
rect 143448 79772 143500 79824
rect 143678 79772 143730 79824
rect 143264 79636 143316 79688
rect 143540 79636 143592 79688
rect 142712 79568 142764 79620
rect 142896 79568 142948 79620
rect 143954 79772 144006 79824
rect 144092 79704 144144 79756
rect 143908 79636 143960 79688
rect 144782 79772 144834 79824
rect 144920 79704 144972 79756
rect 145012 79704 145064 79756
rect 144276 79568 144328 79620
rect 144736 79568 144788 79620
rect 144828 79568 144880 79620
rect 144000 79500 144052 79552
rect 144552 79500 144604 79552
rect 145012 79500 145064 79552
rect 145426 79772 145478 79824
rect 145610 79908 145662 79960
rect 145702 79908 145754 79960
rect 145656 79772 145708 79824
rect 145886 79908 145938 79960
rect 146162 79908 146214 79960
rect 146438 79908 146490 79960
rect 146622 79908 146674 79960
rect 146714 79908 146766 79960
rect 147174 79908 147226 79960
rect 147266 79908 147318 79960
rect 147450 79908 147502 79960
rect 147910 79908 147962 79960
rect 148278 79908 148330 79960
rect 149198 79908 149250 79960
rect 149842 79908 149894 79960
rect 149934 79908 149986 79960
rect 150026 79908 150078 79960
rect 150118 79908 150170 79960
rect 145978 79840 146030 79892
rect 145932 79704 145984 79756
rect 146024 79636 146076 79688
rect 145380 79568 145432 79620
rect 145472 79568 145524 79620
rect 145748 79568 145800 79620
rect 146484 79568 146536 79620
rect 146392 79500 146444 79552
rect 146898 79840 146950 79892
rect 146852 79636 146904 79688
rect 147082 79840 147134 79892
rect 147312 79772 147364 79824
rect 147634 79840 147686 79892
rect 147220 79636 147272 79688
rect 147496 79636 147548 79688
rect 146760 79568 146812 79620
rect 146944 79568 146996 79620
rect 142620 79432 142672 79484
rect 143816 79432 143868 79484
rect 148922 79840 148974 79892
rect 148186 79772 148238 79824
rect 148324 79772 148376 79824
rect 148232 79636 148284 79688
rect 148692 79500 148744 79552
rect 149290 79772 149342 79824
rect 149244 79568 149296 79620
rect 149152 79500 149204 79552
rect 149336 79500 149388 79552
rect 149658 79840 149710 79892
rect 149888 79704 149940 79756
rect 149980 79704 150032 79756
rect 150072 79704 150124 79756
rect 149796 79636 149848 79688
rect 150164 79568 150216 79620
rect 150486 79908 150538 79960
rect 150578 79908 150630 79960
rect 150762 79908 150814 79960
rect 150946 79908 150998 79960
rect 151038 79840 151090 79892
rect 150808 79772 150860 79824
rect 150900 79704 150952 79756
rect 150716 79636 150768 79688
rect 150992 79568 151044 79620
rect 151406 79908 151458 79960
rect 151314 79840 151366 79892
rect 151452 79704 151504 79756
rect 152142 79908 152194 79960
rect 152234 79840 152286 79892
rect 152004 79568 152056 79620
rect 152418 79908 152470 79960
rect 177028 80316 177080 80368
rect 580540 80656 580592 80708
rect 153246 79908 153298 79960
rect 153706 79908 153758 79960
rect 153890 79908 153942 79960
rect 154258 79908 154310 79960
rect 154626 79908 154678 79960
rect 155822 79908 155874 79960
rect 155914 79908 155966 79960
rect 156006 79908 156058 79960
rect 156098 79908 156150 79960
rect 156466 79908 156518 79960
rect 156742 79908 156794 79960
rect 156926 79908 156978 79960
rect 157018 79908 157070 79960
rect 157202 79908 157254 79960
rect 153430 79840 153482 79892
rect 152786 79772 152838 79824
rect 153200 79772 153252 79824
rect 152740 79636 152792 79688
rect 153384 79636 153436 79688
rect 150440 79500 150492 79552
rect 151268 79500 151320 79552
rect 151820 79500 151872 79552
rect 152280 79500 152332 79552
rect 153798 79840 153850 79892
rect 154166 79840 154218 79892
rect 153752 79704 153804 79756
rect 153844 79704 153896 79756
rect 154902 79840 154954 79892
rect 155178 79840 155230 79892
rect 155454 79840 155506 79892
rect 154212 79704 154264 79756
rect 154488 79636 154540 79688
rect 154580 79636 154632 79688
rect 154764 79568 154816 79620
rect 155408 79704 155460 79756
rect 155776 79704 155828 79756
rect 155868 79704 155920 79756
rect 155316 79568 155368 79620
rect 154028 79500 154080 79552
rect 155500 79500 155552 79552
rect 156282 79840 156334 79892
rect 156558 79840 156610 79892
rect 156650 79840 156702 79892
rect 156328 79636 156380 79688
rect 156420 79636 156472 79688
rect 156512 79636 156564 79688
rect 156696 79636 156748 79688
rect 156788 79636 156840 79688
rect 156052 79568 156104 79620
rect 156236 79500 156288 79552
rect 157156 79772 157208 79824
rect 157064 79568 157116 79620
rect 157156 79500 157208 79552
rect 157248 79500 157300 79552
rect 157754 79908 157806 79960
rect 158398 79908 158450 79960
rect 158674 79908 158726 79960
rect 158766 79908 158818 79960
rect 159134 79908 159186 79960
rect 159870 79908 159922 79960
rect 159962 79908 160014 79960
rect 160146 79908 160198 79960
rect 160514 79908 160566 79960
rect 160606 79908 160658 79960
rect 160974 79908 161026 79960
rect 157478 79840 157530 79892
rect 157662 79840 157714 79892
rect 157846 79840 157898 79892
rect 157616 79568 157668 79620
rect 158214 79772 158266 79824
rect 158490 79840 158542 79892
rect 158444 79704 158496 79756
rect 158168 79636 158220 79688
rect 157892 79568 157944 79620
rect 158352 79568 158404 79620
rect 158858 79840 158910 79892
rect 158812 79704 158864 79756
rect 159042 79840 159094 79892
rect 159226 79840 159278 79892
rect 159410 79840 159462 79892
rect 159364 79704 159416 79756
rect 159088 79636 159140 79688
rect 159180 79636 159232 79688
rect 158996 79568 159048 79620
rect 159594 79840 159646 79892
rect 159548 79704 159600 79756
rect 160054 79840 160106 79892
rect 160008 79568 160060 79620
rect 160192 79568 160244 79620
rect 157524 79500 157576 79552
rect 157708 79500 157760 79552
rect 159640 79500 159692 79552
rect 159824 79500 159876 79552
rect 160100 79500 160152 79552
rect 160376 79500 160428 79552
rect 160698 79772 160750 79824
rect 160928 79772 160980 79824
rect 161250 79908 161302 79960
rect 161526 79908 161578 79960
rect 161802 79908 161854 79960
rect 161158 79840 161210 79892
rect 161342 79772 161394 79824
rect 160928 79636 160980 79688
rect 161112 79636 161164 79688
rect 161572 79704 161624 79756
rect 161388 79636 161440 79688
rect 161020 79568 161072 79620
rect 161296 79568 161348 79620
rect 147956 79432 148008 79484
rect 148324 79432 148376 79484
rect 127900 79296 127952 79348
rect 128728 79296 128780 79348
rect 143080 79364 143132 79416
rect 143540 79364 143592 79416
rect 161756 79432 161808 79484
rect 162262 79908 162314 79960
rect 162446 79908 162498 79960
rect 162538 79908 162590 79960
rect 162814 79908 162866 79960
rect 162078 79772 162130 79824
rect 162170 79772 162222 79824
rect 162354 79772 162406 79824
rect 162446 79772 162498 79824
rect 162124 79636 162176 79688
rect 162216 79636 162268 79688
rect 162308 79636 162360 79688
rect 162630 79772 162682 79824
rect 162676 79636 162728 79688
rect 162492 79568 162544 79620
rect 162584 79500 162636 79552
rect 163090 79908 163142 79960
rect 163458 79908 163510 79960
rect 163642 79908 163694 79960
rect 163918 79908 163970 79960
rect 164010 79908 164062 79960
rect 162952 79636 163004 79688
rect 162952 79500 163004 79552
rect 163504 79500 163556 79552
rect 162676 79432 162728 79484
rect 163136 79432 163188 79484
rect 163826 79772 163878 79824
rect 163964 79636 164016 79688
rect 164056 79636 164108 79688
rect 163872 79568 163924 79620
rect 163780 79432 163832 79484
rect 164286 79908 164338 79960
rect 164654 79908 164706 79960
rect 164838 79908 164890 79960
rect 164930 79908 164982 79960
rect 164470 79840 164522 79892
rect 164240 79636 164292 79688
rect 164608 79568 164660 79620
rect 164700 79500 164752 79552
rect 164516 79432 164568 79484
rect 165574 79908 165626 79960
rect 165666 79908 165718 79960
rect 165942 79908 165994 79960
rect 166310 79908 166362 79960
rect 165298 79840 165350 79892
rect 164976 79772 165028 79824
rect 165206 79772 165258 79824
rect 165068 79704 165120 79756
rect 164976 79636 165028 79688
rect 165758 79772 165810 79824
rect 165988 79772 166040 79824
rect 165896 79704 165948 79756
rect 165344 79568 165396 79620
rect 165620 79568 165672 79620
rect 165896 79568 165948 79620
rect 165252 79500 165304 79552
rect 165804 79500 165856 79552
rect 165160 79432 165212 79484
rect 165436 79432 165488 79484
rect 166586 79908 166638 79960
rect 166678 79908 166730 79960
rect 166770 79908 166822 79960
rect 166862 79908 166914 79960
rect 166632 79704 166684 79756
rect 166540 79568 166592 79620
rect 166908 79704 166960 79756
rect 167414 79908 167466 79960
rect 167506 79908 167558 79960
rect 167598 79908 167650 79960
rect 167690 79908 167742 79960
rect 167782 79908 167834 79960
rect 167966 79908 168018 79960
rect 167230 79840 167282 79892
rect 167460 79636 167512 79688
rect 167276 79568 167328 79620
rect 167368 79568 167420 79620
rect 167874 79840 167926 79892
rect 167644 79704 167696 79756
rect 167736 79704 167788 79756
rect 167828 79568 167880 79620
rect 166908 79500 166960 79552
rect 167000 79500 167052 79552
rect 167460 79500 167512 79552
rect 166724 79432 166776 79484
rect 167184 79432 167236 79484
rect 168334 79908 168386 79960
rect 168426 79908 168478 79960
rect 168150 79840 168202 79892
rect 168288 79772 168340 79824
rect 168380 79772 168432 79824
rect 168104 79636 168156 79688
rect 168196 79636 168248 79688
rect 168886 79908 168938 79960
rect 169070 79908 169122 79960
rect 168702 79840 168754 79892
rect 169162 79840 169214 79892
rect 168932 79772 168984 79824
rect 169024 79772 169076 79824
rect 169254 79772 169306 79824
rect 169346 79772 169398 79824
rect 169116 79704 169168 79756
rect 168840 79568 168892 79620
rect 168380 79500 168432 79552
rect 169208 79568 169260 79620
rect 169530 79908 169582 79960
rect 169990 79908 170042 79960
rect 170082 79908 170134 79960
rect 170174 79908 170226 79960
rect 170358 79908 170410 79960
rect 170542 79908 170594 79960
rect 170634 79908 170686 79960
rect 169622 79840 169674 79892
rect 169714 79840 169766 79892
rect 169806 79840 169858 79892
rect 169576 79704 169628 79756
rect 169668 79704 169720 79756
rect 169944 79772 169996 79824
rect 169760 79636 169812 79688
rect 169484 79568 169536 79620
rect 170036 79636 170088 79688
rect 170496 79772 170548 79824
rect 174452 80248 174504 80300
rect 180156 80248 180208 80300
rect 171186 79908 171238 79960
rect 170404 79704 170456 79756
rect 170588 79704 170640 79756
rect 170128 79568 170180 79620
rect 171738 79840 171790 79892
rect 172014 79908 172066 79960
rect 174452 80112 174504 80164
rect 178592 80180 178644 80232
rect 356060 80180 356112 80232
rect 374000 80112 374052 80164
rect 174544 80044 174596 80096
rect 426440 80044 426492 80096
rect 175280 79976 175332 80028
rect 173118 79908 173170 79960
rect 173210 79908 173262 79960
rect 172934 79840 172986 79892
rect 173072 79772 173124 79824
rect 172980 79704 173032 79756
rect 173486 79908 173538 79960
rect 173578 79908 173630 79960
rect 173762 79908 173814 79960
rect 173854 79908 173906 79960
rect 174038 79908 174090 79960
rect 174360 79908 174412 79960
rect 173394 79840 173446 79892
rect 173348 79704 173400 79756
rect 173532 79704 173584 79756
rect 173900 79772 173952 79824
rect 171600 79636 171652 79688
rect 173164 79636 173216 79688
rect 173900 79636 173952 79688
rect 173992 79636 174044 79688
rect 171508 79568 171560 79620
rect 172060 79568 172112 79620
rect 172520 79568 172572 79620
rect 169852 79500 169904 79552
rect 170312 79500 170364 79552
rect 171600 79500 171652 79552
rect 176292 79568 176344 79620
rect 172704 79500 172756 79552
rect 173072 79500 173124 79552
rect 173716 79500 173768 79552
rect 171324 79432 171376 79484
rect 171784 79432 171836 79484
rect 177028 79432 177080 79484
rect 152556 79296 152608 79348
rect 153108 79296 153160 79348
rect 160744 79296 160796 79348
rect 171140 79296 171192 79348
rect 180248 79364 180300 79416
rect 527180 79364 527232 79416
rect 171968 79296 172020 79348
rect 172520 79296 172572 79348
rect 580080 79296 580132 79348
rect 120632 79228 120684 79280
rect 167000 79228 167052 79280
rect 168012 79228 168064 79280
rect 173900 79228 173952 79280
rect 128728 79092 128780 79144
rect 143540 79160 143592 79212
rect 153200 79160 153252 79212
rect 157708 79160 157760 79212
rect 160376 79160 160428 79212
rect 160560 79160 160612 79212
rect 160744 79160 160796 79212
rect 171324 79160 171376 79212
rect 173992 79160 174044 79212
rect 127900 79024 127952 79076
rect 137100 79024 137152 79076
rect 152648 79024 152700 79076
rect 153016 79024 153068 79076
rect 154580 79024 154632 79076
rect 172336 79092 172388 79144
rect 172428 79092 172480 79144
rect 175924 79092 175976 79144
rect 171692 79024 171744 79076
rect 398196 79024 398248 79076
rect 159180 78956 159232 79008
rect 430580 78956 430632 79008
rect 127440 78888 127492 78940
rect 127716 78888 127768 78940
rect 137100 78888 137152 78940
rect 148324 78888 148376 78940
rect 151912 78888 151964 78940
rect 152648 78888 152700 78940
rect 157800 78888 157852 78940
rect 164056 78888 164108 78940
rect 125968 78820 126020 78872
rect 127532 78820 127584 78872
rect 152556 78820 152608 78872
rect 163136 78820 163188 78872
rect 127716 78752 127768 78804
rect 129372 78752 129424 78804
rect 152096 78752 152148 78804
rect 154396 78752 154448 78804
rect 154948 78752 155000 78804
rect 155132 78752 155184 78804
rect 156420 78752 156472 78804
rect 160376 78752 160428 78804
rect 161572 78752 161624 78804
rect 171416 78888 171468 78940
rect 172060 78888 172112 78940
rect 173256 78888 173308 78940
rect 176108 78888 176160 78940
rect 504364 78888 504416 78940
rect 165712 78820 165764 78872
rect 166172 78820 166224 78872
rect 167460 78820 167512 78872
rect 532700 78820 532752 78872
rect 168472 78752 168524 78804
rect 168656 78752 168708 78804
rect 168932 78752 168984 78804
rect 554780 78752 554832 78804
rect 151452 78684 151504 78736
rect 153200 78684 153252 78736
rect 164240 78684 164292 78736
rect 169576 78684 169628 78736
rect 170312 78684 170364 78736
rect 557540 78684 557592 78736
rect 128360 78616 128412 78668
rect 131580 78616 131632 78668
rect 135536 78616 135588 78668
rect 135904 78616 135956 78668
rect 136824 78616 136876 78668
rect 137376 78616 137428 78668
rect 138112 78616 138164 78668
rect 138572 78616 138624 78668
rect 140872 78616 140924 78668
rect 141516 78616 141568 78668
rect 153384 78616 153436 78668
rect 153660 78616 153712 78668
rect 160928 78616 160980 78668
rect 162400 78616 162452 78668
rect 164424 78616 164476 78668
rect 164608 78616 164660 78668
rect 122196 78412 122248 78464
rect 128544 78548 128596 78600
rect 137008 78548 137060 78600
rect 137192 78548 137244 78600
rect 138940 78548 138992 78600
rect 139124 78548 139176 78600
rect 150440 78548 150492 78600
rect 156972 78548 157024 78600
rect 159640 78548 159692 78600
rect 168012 78548 168064 78600
rect 128544 78412 128596 78464
rect 132868 78412 132920 78464
rect 147680 78412 147732 78464
rect 164608 78480 164660 78532
rect 166172 78480 166224 78532
rect 166356 78480 166408 78532
rect 167000 78480 167052 78532
rect 174176 78548 174228 78600
rect 175648 78548 175700 78600
rect 398104 78616 398156 78668
rect 172152 78480 172204 78532
rect 180064 78480 180116 78532
rect 160376 78412 160428 78464
rect 172060 78412 172112 78464
rect 173256 78412 173308 78464
rect 397552 78480 397604 78532
rect 116584 78344 116636 78396
rect 129188 78344 129240 78396
rect 141056 78344 141108 78396
rect 171600 78344 171652 78396
rect 171876 78344 171928 78396
rect 179972 78344 180024 78396
rect 114560 78276 114612 78328
rect 134432 78276 134484 78328
rect 138388 78276 138440 78328
rect 138756 78276 138808 78328
rect 139952 78276 140004 78328
rect 178040 78276 178092 78328
rect 113824 78208 113876 78260
rect 125324 78208 125376 78260
rect 131580 78208 131632 78260
rect 132132 78208 132184 78260
rect 134064 78208 134116 78260
rect 134248 78208 134300 78260
rect 141056 78208 141108 78260
rect 141608 78208 141660 78260
rect 161572 78208 161624 78260
rect 162124 78208 162176 78260
rect 162400 78208 162452 78260
rect 242164 78208 242216 78260
rect 110420 78140 110472 78192
rect 122932 78140 122984 78192
rect 123300 78140 123352 78192
rect 107660 78072 107712 78124
rect 123392 78072 123444 78124
rect 126060 78140 126112 78192
rect 126336 78140 126388 78192
rect 126428 78140 126480 78192
rect 130476 78140 130528 78192
rect 133880 78140 133932 78192
rect 135996 78140 136048 78192
rect 144184 78140 144236 78192
rect 152556 78140 152608 78192
rect 159364 78140 159416 78192
rect 162952 78140 163004 78192
rect 93124 78004 93176 78056
rect 125968 78004 126020 78056
rect 127900 78072 127952 78124
rect 135444 78072 135496 78124
rect 132776 78004 132828 78056
rect 134248 78004 134300 78056
rect 134892 78004 134944 78056
rect 135996 78004 136048 78056
rect 136180 78004 136232 78056
rect 89720 77936 89772 77988
rect 123300 77936 123352 77988
rect 124956 77936 125008 77988
rect 127072 77936 127124 77988
rect 127440 77936 127492 77988
rect 127624 77936 127676 77988
rect 130200 77936 130252 77988
rect 130384 77936 130436 77988
rect 131304 77936 131356 77988
rect 132040 77936 132092 77988
rect 134432 77936 134484 77988
rect 134800 77936 134852 77988
rect 139676 77936 139728 77988
rect 160928 78072 160980 78124
rect 161664 78072 161716 78124
rect 304264 78140 304316 78192
rect 157064 78004 157116 78056
rect 155500 77936 155552 77988
rect 159640 77936 159692 77988
rect 162952 77936 163004 77988
rect 169392 77936 169444 77988
rect 125324 77868 125376 77920
rect 133420 77868 133472 77920
rect 142068 77868 142120 77920
rect 152188 77868 152240 77920
rect 120080 77800 120132 77852
rect 124036 77800 124088 77852
rect 124128 77800 124180 77852
rect 135352 77800 135404 77852
rect 144920 77800 144972 77852
rect 164240 77868 164292 77920
rect 169576 78072 169628 78124
rect 498200 78072 498252 78124
rect 170588 78004 170640 78056
rect 574744 78004 574796 78056
rect 170772 77936 170824 77988
rect 581092 77936 581144 77988
rect 171968 77868 172020 77920
rect 172060 77868 172112 77920
rect 173624 77868 173676 77920
rect 173992 77868 174044 77920
rect 174452 77868 174504 77920
rect 152556 77800 152608 77852
rect 162124 77800 162176 77852
rect 165896 77800 165948 77852
rect 170588 77800 170640 77852
rect 171324 77800 171376 77852
rect 172428 77800 172480 77852
rect 129188 77732 129240 77784
rect 129832 77732 129884 77784
rect 131304 77732 131356 77784
rect 131764 77732 131816 77784
rect 159180 77732 159232 77784
rect 158904 77664 158956 77716
rect 164056 77732 164108 77784
rect 172244 77732 172296 77784
rect 125140 77596 125192 77648
rect 126704 77596 126756 77648
rect 155868 77596 155920 77648
rect 162492 77596 162544 77648
rect 171784 77664 171836 77716
rect 171692 77596 171744 77648
rect 123392 77528 123444 77580
rect 129740 77528 129792 77580
rect 147680 77528 147732 77580
rect 148048 77528 148100 77580
rect 154672 77528 154724 77580
rect 158260 77528 158312 77580
rect 159916 77528 159968 77580
rect 172060 77528 172112 77580
rect 122932 77460 122984 77512
rect 134064 77460 134116 77512
rect 152188 77460 152240 77512
rect 152832 77460 152884 77512
rect 154488 77460 154540 77512
rect 158628 77460 158680 77512
rect 163136 77460 163188 77512
rect 173348 77460 173400 77512
rect 123576 77392 123628 77444
rect 134984 77392 135036 77444
rect 154028 77392 154080 77444
rect 120816 77324 120868 77376
rect 128084 77324 128136 77376
rect 150348 77324 150400 77376
rect 153108 77324 153160 77376
rect 153384 77324 153436 77376
rect 154120 77324 154172 77376
rect 154672 77392 154724 77444
rect 155316 77392 155368 77444
rect 157432 77392 157484 77444
rect 157984 77392 158036 77444
rect 169392 77392 169444 77444
rect 175924 77392 175976 77444
rect 180064 77392 180116 77444
rect 396724 77392 396776 77444
rect 155224 77324 155276 77376
rect 155408 77324 155460 77376
rect 155684 77324 155736 77376
rect 127072 77256 127124 77308
rect 127900 77256 127952 77308
rect 130476 77256 130528 77308
rect 135812 77256 135864 77308
rect 149520 77256 149572 77308
rect 149704 77256 149756 77308
rect 152188 77256 152240 77308
rect 152464 77256 152516 77308
rect 154212 77256 154264 77308
rect 155500 77256 155552 77308
rect 156420 77256 156472 77308
rect 156696 77256 156748 77308
rect 119436 77188 119488 77240
rect 172888 77188 172940 77240
rect 143172 77120 143224 77172
rect 226340 77120 226392 77172
rect 123484 76984 123536 77036
rect 132316 76984 132368 77036
rect 147956 76984 148008 77036
rect 148416 76984 148468 77036
rect 149244 76984 149296 77036
rect 149980 76984 150032 77036
rect 124864 76916 124916 76968
rect 135168 76916 135220 76968
rect 149152 76916 149204 76968
rect 149612 76916 149664 76968
rect 150164 76916 150216 76968
rect 168840 77052 168892 77104
rect 171784 77052 171836 77104
rect 249800 77052 249852 77104
rect 118700 76848 118752 76900
rect 134616 76848 134668 76900
rect 144828 76848 144880 76900
rect 247040 76984 247092 77036
rect 168840 76916 168892 76968
rect 260840 76916 260892 76968
rect 164608 76848 164660 76900
rect 284300 76848 284352 76900
rect 102140 76780 102192 76832
rect 132684 76780 132736 76832
rect 143724 76780 143776 76832
rect 144368 76780 144420 76832
rect 148600 76780 148652 76832
rect 296720 76780 296772 76832
rect 70400 76712 70452 76764
rect 131212 76712 131264 76764
rect 135168 76712 135220 76764
rect 138020 76712 138072 76764
rect 148048 76712 148100 76764
rect 148324 76712 148376 76764
rect 149244 76712 149296 76764
rect 149888 76712 149940 76764
rect 152280 76712 152332 76764
rect 152740 76712 152792 76764
rect 157616 76712 157668 76764
rect 157892 76712 157944 76764
rect 164240 76712 164292 76764
rect 171784 76712 171836 76764
rect 172336 76712 172388 76764
rect 376760 76712 376812 76764
rect 93860 76644 93912 76696
rect 128544 76644 128596 76696
rect 137928 76644 137980 76696
rect 144368 76644 144420 76696
rect 147864 76644 147916 76696
rect 148232 76644 148284 76696
rect 154856 76644 154908 76696
rect 375380 76644 375432 76696
rect 69020 76576 69072 76628
rect 130936 76576 130988 76628
rect 157616 76576 157668 76628
rect 158076 76576 158128 76628
rect 160100 76576 160152 76628
rect 444380 76576 444432 76628
rect 6920 76508 6972 76560
rect 124772 76508 124824 76560
rect 147680 76508 147732 76560
rect 147864 76508 147916 76560
rect 154856 76508 154908 76560
rect 155408 76508 155460 76560
rect 165620 76508 165672 76560
rect 170680 76508 170732 76560
rect 171600 76508 171652 76560
rect 171876 76508 171928 76560
rect 132960 76440 133012 76492
rect 133236 76440 133288 76492
rect 140412 76440 140464 76492
rect 147680 76372 147732 76424
rect 148508 76372 148560 76424
rect 139308 76304 139360 76356
rect 140412 76304 140464 76356
rect 147036 76236 147088 76288
rect 168564 76440 168616 76492
rect 168932 76440 168984 76492
rect 169024 76440 169076 76492
rect 558920 76508 558972 76560
rect 170956 76372 171008 76424
rect 173348 76372 173400 76424
rect 171416 76304 171468 76356
rect 172336 76304 172388 76356
rect 190460 76440 190512 76492
rect 140780 76032 140832 76084
rect 141148 76032 141200 76084
rect 145012 76032 145064 76084
rect 124036 75964 124088 76016
rect 120724 75896 120776 75948
rect 145104 75964 145156 76016
rect 145380 75964 145432 76016
rect 145656 75964 145708 76016
rect 139676 75896 139728 75948
rect 140044 75896 140096 75948
rect 141148 75896 141200 75948
rect 141700 75896 141752 75948
rect 144184 75896 144236 75948
rect 144736 75896 144788 75948
rect 146852 76168 146904 76220
rect 146668 76100 146720 76152
rect 147036 76100 147088 76152
rect 146484 76032 146536 76084
rect 146852 76032 146904 76084
rect 146668 75964 146720 76016
rect 160100 76168 160152 76220
rect 160560 76168 160612 76220
rect 165804 76168 165856 76220
rect 166816 76168 166868 76220
rect 150440 75964 150492 76016
rect 150624 75964 150676 76016
rect 146484 75896 146536 75948
rect 146576 75896 146628 75948
rect 147220 75896 147272 75948
rect 158904 75896 158956 75948
rect 159456 75896 159508 75948
rect 160652 76100 160704 76152
rect 161756 76100 161808 76152
rect 161940 76100 161992 76152
rect 163412 76100 163464 76152
rect 162860 76032 162912 76084
rect 162952 76032 163004 76084
rect 163964 76032 164016 76084
rect 161756 75964 161808 76016
rect 162032 75964 162084 76016
rect 163136 75964 163188 76016
rect 163872 75964 163924 76016
rect 160560 75896 160612 75948
rect 161480 75896 161532 75948
rect 162216 75896 162268 75948
rect 163412 75896 163464 75948
rect 163688 75896 163740 75948
rect 164608 75896 164660 75948
rect 165252 75896 165304 75948
rect 165436 75896 165488 75948
rect 165804 75896 165856 75948
rect 165896 75896 165948 75948
rect 166632 75896 166684 75948
rect 166908 75896 166960 75948
rect 167368 75896 167420 75948
rect 167460 75896 167512 75948
rect 167736 75896 167788 75948
rect 172704 75828 172756 75880
rect 172520 75760 172572 75812
rect 139952 75692 140004 75744
rect 140228 75692 140280 75744
rect 159088 75692 159140 75744
rect 159824 75692 159876 75744
rect 160100 75692 160152 75744
rect 161020 75692 161072 75744
rect 167368 75692 167420 75744
rect 167644 75692 167696 75744
rect 139584 75624 139636 75676
rect 140136 75624 140188 75676
rect 157340 75624 157392 75676
rect 158168 75624 158220 75676
rect 75920 75420 75972 75472
rect 132040 75556 132092 75608
rect 121460 75488 121512 75540
rect 134616 75488 134668 75540
rect 162584 75488 162636 75540
rect 127164 75420 127216 75472
rect 127716 75420 127768 75472
rect 159732 75420 159784 75472
rect 169944 75488 169996 75540
rect 170312 75488 170364 75540
rect 51080 75352 51132 75404
rect 129004 75352 129056 75404
rect 137100 75352 137152 75404
rect 137744 75352 137796 75404
rect 150808 75352 150860 75404
rect 163780 75352 163832 75404
rect 431960 75420 432012 75472
rect 438860 75352 438912 75404
rect 49700 75284 49752 75336
rect 127164 75284 127216 75336
rect 127256 75284 127308 75336
rect 128084 75284 128136 75336
rect 128544 75284 128596 75336
rect 129648 75284 129700 75336
rect 132684 75284 132736 75336
rect 133604 75284 133656 75336
rect 135352 75284 135404 75336
rect 135628 75284 135680 75336
rect 135812 75284 135864 75336
rect 136456 75284 136508 75336
rect 164884 75284 164936 75336
rect 481640 75284 481692 75336
rect 46940 75216 46992 75268
rect 26240 75148 26292 75200
rect 125968 75148 126020 75200
rect 126888 75148 126940 75200
rect 127164 75148 127216 75200
rect 127808 75148 127860 75200
rect 127072 75080 127124 75132
rect 127440 75080 127492 75132
rect 128728 75216 128780 75268
rect 129096 75216 129148 75268
rect 130016 75216 130068 75268
rect 130660 75216 130712 75268
rect 131396 75216 131448 75268
rect 131948 75216 132000 75268
rect 133052 75216 133104 75268
rect 133788 75216 133840 75268
rect 134156 75216 134208 75268
rect 134524 75216 134576 75268
rect 135720 75216 135772 75268
rect 136272 75216 136324 75268
rect 137100 75216 137152 75268
rect 137468 75216 137520 75268
rect 138296 75216 138348 75268
rect 138480 75216 138532 75268
rect 150808 75216 150860 75268
rect 151176 75216 151228 75268
rect 153200 75216 153252 75268
rect 154120 75216 154172 75268
rect 163872 75216 163924 75268
rect 489920 75216 489972 75268
rect 128636 75148 128688 75200
rect 129556 75148 129608 75200
rect 129740 75148 129792 75200
rect 130476 75148 130528 75200
rect 131212 75148 131264 75200
rect 132132 75148 132184 75200
rect 132776 75148 132828 75200
rect 133696 75148 133748 75200
rect 135628 75148 135680 75200
rect 135996 75148 136048 75200
rect 150624 75148 150676 75200
rect 151084 75148 151136 75200
rect 156236 75148 156288 75200
rect 156512 75148 156564 75200
rect 169760 75148 169812 75200
rect 170036 75148 170088 75200
rect 129372 75080 129424 75132
rect 135444 75080 135496 75132
rect 136364 75080 136416 75132
rect 138296 75080 138348 75132
rect 138572 75080 138624 75132
rect 151912 75080 151964 75132
rect 152464 75080 152516 75132
rect 168840 75080 168892 75132
rect 169208 75080 169260 75132
rect 127992 75012 128044 75064
rect 156052 75012 156104 75064
rect 156512 75012 156564 75064
rect 169760 75012 169812 75064
rect 170220 75012 170272 75064
rect 127440 74944 127492 74996
rect 128268 74944 128320 74996
rect 151912 74944 151964 74996
rect 153016 74944 153068 74996
rect 158812 74944 158864 74996
rect 159272 74944 159324 74996
rect 169300 74944 169352 74996
rect 564440 75148 564492 75200
rect 156052 74876 156104 74928
rect 156788 74876 156840 74928
rect 130476 74468 130528 74520
rect 135260 74468 135312 74520
rect 138756 74468 138808 74520
rect 140136 74468 140188 74520
rect 142252 74128 142304 74180
rect 142804 74128 142856 74180
rect 4160 73992 4212 74044
rect 126336 73992 126388 74044
rect 118792 73924 118844 73976
rect 134432 73924 134484 73976
rect 141884 73924 141936 73976
rect 209780 73924 209832 73976
rect 60740 73856 60792 73908
rect 130200 73856 130252 73908
rect 147312 73856 147364 73908
rect 223580 73856 223632 73908
rect 153200 73788 153252 73840
rect 318800 73788 318852 73840
rect 145012 73720 145064 73772
rect 145840 73720 145892 73772
rect 137560 73516 137612 73568
rect 142988 73516 143040 73568
rect 161664 73448 161716 73500
rect 162308 73448 162360 73500
rect 126244 73176 126296 73228
rect 130844 73176 130896 73228
rect 171048 73108 171100 73160
rect 580172 73108 580224 73160
rect 145472 72904 145524 72956
rect 145932 72904 145984 72956
rect 149980 72768 150032 72820
rect 305000 72768 305052 72820
rect 149704 72700 149756 72752
rect 307760 72700 307812 72752
rect 149796 72632 149848 72684
rect 311900 72632 311952 72684
rect 151360 72564 151412 72616
rect 332600 72564 332652 72616
rect 154488 72496 154540 72548
rect 340880 72496 340932 72548
rect 96620 72428 96672 72480
rect 133144 72428 133196 72480
rect 158628 72428 158680 72480
rect 368480 72428 368532 72480
rect 124772 72360 124824 72412
rect 125416 72360 125468 72412
rect 3424 71680 3476 71732
rect 17316 71680 17368 71732
rect 139124 71476 139176 71528
rect 171140 71476 171192 71528
rect 155132 71408 155184 71460
rect 382280 71408 382332 71460
rect 157984 71340 158036 71392
rect 408500 71340 408552 71392
rect 163412 71272 163464 71324
rect 490012 71272 490064 71324
rect 164976 71204 165028 71256
rect 507860 71204 507912 71256
rect 166540 71136 166592 71188
rect 523040 71136 523092 71188
rect 168012 71068 168064 71120
rect 536840 71068 536892 71120
rect 167920 71000 167972 71052
rect 539600 71000 539652 71052
rect 137284 70456 137336 70508
rect 138756 70388 138808 70440
rect 166356 69708 166408 69760
rect 518900 69708 518952 69760
rect 169484 69640 169536 69692
rect 564532 69640 564584 69692
rect 140044 68416 140096 68468
rect 184940 68416 184992 68468
rect 159272 68348 159324 68400
rect 218704 68348 218756 68400
rect 156972 68280 157024 68332
rect 320180 68280 320232 68332
rect 138572 67532 138624 67584
rect 140044 67532 140096 67584
rect 139952 67056 140004 67108
rect 189080 67056 189132 67108
rect 157892 66988 157944 67040
rect 412640 66988 412692 67040
rect 167644 66920 167696 66972
rect 543740 66920 543792 66972
rect 170220 66852 170272 66904
rect 569960 66852 570012 66904
rect 155684 65628 155736 65680
rect 367100 65628 367152 65680
rect 166264 65560 166316 65612
rect 525800 65560 525852 65612
rect 170128 65492 170180 65544
rect 572720 65492 572772 65544
rect 152464 64472 152516 64524
rect 338120 64472 338172 64524
rect 152556 64404 152608 64456
rect 339500 64404 339552 64456
rect 156696 64336 156748 64388
rect 390560 64336 390612 64388
rect 162032 64268 162084 64320
rect 463700 64268 463752 64320
rect 163412 64200 163464 64252
rect 487160 64200 487212 64252
rect 170036 64132 170088 64184
rect 568580 64132 568632 64184
rect 142804 62976 142856 63028
rect 224960 62976 225012 63028
rect 152372 62908 152424 62960
rect 340972 62908 341024 62960
rect 161940 62840 161992 62892
rect 465080 62840 465132 62892
rect 170496 62772 170548 62824
rect 514760 62772 514812 62824
rect 149612 61412 149664 61464
rect 303620 61412 303672 61464
rect 102232 61344 102284 61396
rect 125324 61344 125376 61396
rect 138480 61344 138532 61396
rect 152464 61344 152516 61396
rect 157800 61344 157852 61396
rect 415400 61344 415452 61396
rect 182916 60664 182968 60716
rect 580172 60664 580224 60716
rect 120080 60188 120132 60240
rect 123576 60188 123628 60240
rect 151084 60188 151136 60240
rect 331220 60188 331272 60240
rect 153752 60120 153804 60172
rect 362960 60120 363012 60172
rect 156604 60052 156656 60104
rect 396080 60052 396132 60104
rect 159180 59984 159232 60036
rect 427820 59984 427872 60036
rect 3056 59304 3108 59356
rect 180892 59304 180944 59356
rect 158352 58692 158404 58744
rect 374092 58692 374144 58744
rect 159088 58624 159140 58676
rect 440240 58624 440292 58676
rect 150992 57264 151044 57316
rect 325700 57264 325752 57316
rect 95240 57196 95292 57248
rect 125232 57196 125284 57248
rect 157708 57196 157760 57248
rect 415492 57196 415544 57248
rect 88340 55836 88392 55888
rect 125048 55836 125100 55888
rect 13820 51688 13872 51740
rect 125140 51688 125192 51740
rect 153660 50396 153712 50448
rect 357440 50396 357492 50448
rect 171692 50328 171744 50380
rect 425060 50328 425112 50380
rect 171784 49036 171836 49088
rect 418160 49036 418212 49088
rect 163320 48968 163372 49020
rect 485780 48968 485832 49020
rect 118240 46860 118292 46912
rect 580172 46860 580224 46912
rect 3424 45500 3476 45552
rect 174084 45500 174136 45552
rect 67640 44956 67692 45008
rect 130200 44956 130252 45008
rect 30380 44888 30432 44940
rect 127532 44888 127584 44940
rect 27620 44820 27672 44872
rect 127624 44820 127676 44872
rect 45560 37884 45612 37936
rect 116584 37884 116636 37936
rect 7564 36524 7616 36576
rect 124220 36524 124272 36576
rect 148416 35368 148468 35420
rect 291200 35368 291252 35420
rect 159732 35300 159784 35352
rect 382372 35300 382424 35352
rect 162492 35232 162544 35284
rect 390652 35232 390704 35284
rect 38660 35164 38712 35216
rect 122196 35164 122248 35216
rect 160744 35164 160796 35216
rect 447140 35164 447192 35216
rect 142712 33804 142764 33856
rect 219440 33804 219492 33856
rect 144276 33736 144328 33788
rect 234620 33736 234672 33788
rect 173348 33056 173400 33108
rect 580172 33056 580224 33108
rect 141424 32852 141476 32904
rect 198740 32852 198792 32904
rect 141516 32784 141568 32836
rect 201500 32784 201552 32836
rect 148232 32716 148284 32768
rect 285680 32716 285732 32768
rect 148324 32648 148376 32700
rect 287060 32648 287112 32700
rect 150900 32580 150952 32632
rect 321560 32580 321612 32632
rect 3424 32512 3476 32564
rect 7656 32512 7708 32564
rect 152188 32512 152240 32564
rect 346400 32512 346452 32564
rect 152280 32444 152332 32496
rect 349160 32444 349212 32496
rect 31760 32376 31812 32428
rect 120816 32376 120868 32428
rect 161848 32376 161900 32428
rect 466460 32376 466512 32428
rect 304264 31152 304316 31204
rect 465172 31152 465224 31204
rect 166172 31084 166224 31136
rect 524420 31084 524472 31136
rect 167552 31016 167604 31068
rect 535460 31016 535512 31068
rect 142620 29928 142672 29980
rect 215300 29928 215352 29980
rect 156512 29860 156564 29912
rect 391940 29860 391992 29912
rect 157524 29792 157576 29844
rect 409880 29792 409932 29844
rect 157616 29724 157668 29776
rect 416780 29724 416832 29776
rect 158996 29656 159048 29708
rect 434720 29656 434772 29708
rect 167460 29588 167512 29640
rect 542360 29588 542412 29640
rect 141332 28568 141384 28620
rect 201592 28568 201644 28620
rect 141240 28500 141292 28552
rect 204260 28500 204312 28552
rect 141148 28432 141200 28484
rect 208400 28432 208452 28484
rect 154120 28364 154172 28416
rect 332692 28364 332744 28416
rect 155040 28296 155092 28348
rect 378140 28296 378192 28348
rect 160652 28228 160704 28280
rect 454040 28228 454092 28280
rect 139768 27276 139820 27328
rect 179420 27276 179472 27328
rect 139860 27208 139912 27260
rect 183560 27208 183612 27260
rect 139676 27140 139728 27192
rect 186320 27140 186372 27192
rect 142528 27072 142580 27124
rect 218060 27072 218112 27124
rect 172244 27004 172296 27056
rect 411260 27004 411312 27056
rect 156420 26936 156472 26988
rect 398840 26936 398892 26988
rect 168932 26868 168984 26920
rect 560300 26868 560352 26920
rect 140320 25916 140372 25968
rect 176752 25916 176804 25968
rect 148140 25848 148192 25900
rect 289820 25848 289872 25900
rect 157432 25780 157484 25832
rect 414020 25780 414072 25832
rect 168748 25712 168800 25764
rect 556160 25712 556212 25764
rect 168840 25644 168892 25696
rect 563060 25644 563112 25696
rect 169852 25576 169904 25628
rect 571340 25576 571392 25628
rect 169944 25508 169996 25560
rect 572812 25508 572864 25560
rect 148048 24488 148100 24540
rect 292580 24488 292632 24540
rect 167092 24420 167144 24472
rect 534080 24420 534132 24472
rect 167276 24352 167328 24404
rect 538220 24352 538272 24404
rect 167368 24284 167420 24336
rect 540980 24284 541032 24336
rect 167184 24216 167236 24268
rect 545120 24216 545172 24268
rect 168656 24148 168708 24200
rect 552020 24148 552072 24200
rect 3332 24080 3384 24132
rect 181076 24080 181128 24132
rect 182824 24080 182876 24132
rect 579620 24080 579672 24132
rect 3424 23128 3476 23180
rect 173992 23128 174044 23180
rect 172152 23060 172204 23112
rect 397460 23060 397512 23112
rect 161756 22992 161808 23044
rect 467840 22992 467892 23044
rect 166080 22924 166132 22976
rect 516140 22924 516192 22976
rect 165988 22856 166040 22908
rect 520280 22856 520332 22908
rect 165896 22788 165948 22840
rect 527180 22788 527232 22840
rect 118332 22720 118384 22772
rect 580264 22720 580316 22772
rect 152096 21632 152148 21684
rect 343640 21632 343692 21684
rect 172060 21564 172112 21616
rect 440332 21564 440384 21616
rect 158904 21496 158956 21548
rect 436100 21496 436152 21548
rect 163228 21428 163280 21480
rect 484400 21428 484452 21480
rect 11060 21360 11112 21412
rect 126152 21360 126204 21412
rect 163136 21360 163188 21412
rect 491300 21360 491352 21412
rect 145472 20612 145524 20664
rect 262220 20612 262272 20664
rect 150808 20544 150860 20596
rect 329840 20544 329892 20596
rect 145656 20476 145708 20528
rect 255320 20476 255372 20528
rect 255964 20476 256016 20528
rect 456892 20476 456944 20528
rect 242164 20408 242216 20460
rect 449900 20408 449952 20460
rect 160284 20340 160336 20392
rect 445760 20340 445812 20392
rect 160468 20272 160520 20324
rect 448520 20272 448572 20324
rect 160192 20204 160244 20256
rect 448612 20204 448664 20256
rect 160100 20136 160152 20188
rect 451280 20136 451332 20188
rect 160560 20068 160612 20120
rect 452660 20068 452712 20120
rect 160376 20000 160428 20052
rect 455420 20000 455472 20052
rect 163044 19932 163096 19984
rect 481732 19932 481784 19984
rect 145564 19864 145616 19916
rect 259460 19864 259512 19916
rect 144184 18844 144236 18896
rect 241520 18844 241572 18896
rect 171968 18776 172020 18828
rect 404360 18776 404412 18828
rect 158812 18708 158864 18760
rect 433340 18708 433392 18760
rect 63500 18640 63552 18692
rect 126336 18640 126388 18692
rect 168472 18640 168524 18692
rect 553400 18640 553452 18692
rect 42800 18572 42852 18624
rect 128820 18572 128872 18624
rect 168564 18572 168616 18624
rect 556252 18572 556304 18624
rect 142436 17824 142488 17876
rect 216680 17824 216732 17876
rect 147128 17756 147180 17808
rect 269120 17756 269172 17808
rect 147036 17688 147088 17740
rect 273260 17688 273312 17740
rect 146944 17620 146996 17672
rect 276020 17620 276072 17672
rect 172428 17552 172480 17604
rect 347780 17552 347832 17604
rect 157340 17484 157392 17536
rect 419540 17484 419592 17536
rect 160008 17416 160060 17468
rect 441620 17416 441672 17468
rect 162952 17348 163004 17400
rect 492680 17348 492732 17400
rect 164792 17280 164844 17332
rect 503720 17280 503772 17332
rect 165528 17212 165580 17264
rect 514852 17212 514904 17264
rect 144092 16192 144144 16244
rect 237656 16192 237708 16244
rect 152004 16124 152056 16176
rect 342904 16124 342956 16176
rect 153568 16056 153620 16108
rect 361120 16056 361172 16108
rect 156328 15988 156380 16040
rect 395344 15988 395396 16040
rect 156236 15920 156288 15972
rect 398932 15920 398984 15972
rect 156144 15852 156196 15904
rect 402520 15852 402572 15904
rect 145288 15104 145340 15156
rect 254216 15104 254268 15156
rect 145380 15036 145432 15088
rect 258264 15036 258316 15088
rect 146852 14968 146904 15020
rect 268384 14968 268436 15020
rect 146760 14900 146812 14952
rect 272432 14900 272484 14952
rect 149520 14832 149572 14884
rect 311440 14832 311492 14884
rect 154948 14764 155000 14816
rect 379520 14764 379572 14816
rect 154764 14696 154816 14748
rect 381176 14696 381228 14748
rect 154672 14628 154724 14680
rect 384304 14628 384356 14680
rect 154856 14560 154908 14612
rect 386696 14560 386748 14612
rect 164700 14492 164752 14544
rect 500592 14492 500644 14544
rect 165804 14424 165856 14476
rect 523776 14424 523828 14476
rect 145196 14356 145248 14408
rect 251272 14356 251324 14408
rect 139584 14288 139636 14340
rect 188528 14288 188580 14340
rect 151912 13404 151964 13456
rect 349252 13404 349304 13456
rect 153292 13336 153344 13388
rect 357532 13336 357584 13388
rect 153476 13268 153528 13320
rect 359464 13268 359516 13320
rect 155592 13200 155644 13252
rect 361856 13200 361908 13252
rect 153384 13132 153436 13184
rect 365812 13132 365864 13184
rect 162860 13064 162912 13116
rect 488816 13064 488868 13116
rect 143908 12384 143960 12436
rect 236552 12384 236604 12436
rect 146668 12316 146720 12368
rect 276112 12316 276164 12368
rect 150716 12248 150768 12300
rect 328000 12248 328052 12300
rect 150624 12180 150676 12232
rect 328736 12180 328788 12232
rect 151820 12112 151872 12164
rect 345296 12112 345348 12164
rect 156052 12044 156104 12096
rect 400864 12044 400916 12096
rect 161664 11976 161716 12028
rect 473452 11976 473504 12028
rect 164332 11908 164384 11960
rect 498936 11908 498988 11960
rect 164424 11840 164476 11892
rect 502984 11840 503036 11892
rect 117320 11772 117372 11824
rect 134248 11772 134300 11824
rect 164516 11772 164568 11824
rect 506480 11772 506532 11824
rect 106464 11704 106516 11756
rect 133052 11704 133104 11756
rect 164608 11704 164660 11756
rect 509608 11704 509660 11756
rect 144000 11636 144052 11688
rect 233424 11636 233476 11688
rect 162400 11568 162452 11620
rect 240140 11568 240192 11620
rect 139492 11500 139544 11552
rect 176660 11432 176712 11484
rect 177856 11432 177908 11484
rect 184940 11500 184992 11552
rect 186136 11500 186188 11552
rect 201500 11500 201552 11552
rect 202696 11500 202748 11552
rect 184940 11364 184992 11416
rect 85672 10548 85724 10600
rect 131672 10548 131724 10600
rect 81624 10480 81676 10532
rect 131764 10480 131816 10532
rect 78128 10412 78180 10464
rect 128360 10412 128412 10464
rect 150532 10412 150584 10464
rect 324412 10412 324464 10464
rect 25320 10344 25372 10396
rect 93124 10344 93176 10396
rect 99840 10344 99892 10396
rect 132960 10344 133012 10396
rect 161572 10344 161624 10396
rect 469864 10344 469916 10396
rect 35992 10276 36044 10328
rect 127440 10276 127492 10328
rect 167000 10276 167052 10328
rect 539692 10276 539744 10328
rect 146576 9528 146628 9580
rect 278320 9528 278372 9580
rect 147864 9460 147916 9512
rect 288992 9460 289044 9512
rect 147956 9392 148008 9444
rect 292580 9392 292632 9444
rect 147772 9324 147824 9376
rect 296076 9324 296128 9376
rect 60832 9256 60884 9308
rect 129004 9256 129056 9308
rect 149152 9256 149204 9308
rect 303160 9256 303212 9308
rect 59636 9188 59688 9240
rect 130108 9188 130160 9240
rect 149428 9188 149480 9240
rect 306748 9188 306800 9240
rect 52552 9120 52604 9172
rect 128636 9120 128688 9172
rect 149336 9120 149388 9172
rect 310244 9120 310296 9172
rect 53748 9052 53800 9104
rect 128544 9052 128596 9104
rect 149244 9052 149296 9104
rect 313832 9052 313884 9104
rect 45468 8984 45520 9036
rect 128728 8984 128780 9036
rect 165436 8984 165488 9036
rect 507676 8984 507728 9036
rect 9956 8916 10008 8968
rect 126060 8916 126112 8968
rect 165712 8916 165764 8968
rect 521844 8916 521896 8968
rect 116400 7964 116452 8016
rect 134156 7964 134208 8016
rect 105728 7896 105780 7948
rect 132776 7896 132828 7948
rect 98644 7828 98696 7880
rect 132868 7828 132920 7880
rect 142252 7828 142304 7880
rect 222752 7828 222804 7880
rect 84476 7760 84528 7812
rect 131580 7760 131632 7812
rect 149060 7760 149112 7812
rect 307944 7760 307996 7812
rect 48964 7692 49016 7744
rect 129188 7692 129240 7744
rect 150440 7692 150492 7744
rect 323308 7692 323360 7744
rect 34796 7624 34848 7676
rect 127348 7624 127400 7676
rect 155868 7624 155920 7676
rect 385960 7624 386012 7676
rect 24216 7556 24268 7608
rect 122104 7556 122156 7608
rect 158720 7556 158772 7608
rect 429660 7556 429712 7608
rect 139400 6808 139452 6860
rect 181444 6808 181496 6860
rect 143816 6740 143868 6792
rect 239312 6740 239364 6792
rect 143724 6672 143776 6724
rect 242992 6672 243044 6724
rect 104532 6604 104584 6656
rect 132684 6604 132736 6656
rect 145104 6604 145156 6656
rect 253480 6604 253532 6656
rect 80888 6536 80940 6588
rect 131396 6536 131448 6588
rect 144920 6536 144972 6588
rect 257068 6536 257120 6588
rect 77392 6468 77444 6520
rect 131488 6468 131540 6520
rect 145012 6468 145064 6520
rect 260656 6468 260708 6520
rect 66720 6400 66772 6452
rect 130016 6400 130068 6452
rect 146392 6400 146444 6452
rect 271236 6400 271288 6452
rect 44272 6332 44324 6384
rect 128912 6332 128964 6384
rect 146484 6332 146536 6384
rect 274824 6332 274876 6384
rect 33600 6264 33652 6316
rect 127256 6264 127308 6316
rect 137008 6264 137060 6316
rect 149520 6264 149572 6316
rect 155960 6264 156012 6316
rect 394240 6264 394292 6316
rect 19432 6196 19484 6248
rect 124956 6196 125008 6248
rect 137100 6196 137152 6248
rect 154212 6196 154264 6248
rect 161480 6196 161532 6248
rect 471060 6196 471112 6248
rect 18236 6128 18288 6180
rect 125968 6128 126020 6180
rect 137192 6128 137244 6180
rect 157800 6128 157852 6180
rect 168380 6128 168432 6180
rect 562048 6128 562100 6180
rect 108304 5312 108356 5364
rect 113824 5312 113876 5364
rect 114008 5312 114060 5364
rect 134064 5312 134116 5364
rect 101036 5244 101088 5296
rect 133144 5244 133196 5296
rect 93952 5176 94004 5228
rect 133328 5176 133380 5228
rect 138112 5176 138164 5228
rect 166080 5176 166132 5228
rect 63224 5108 63276 5160
rect 129924 5108 129976 5160
rect 141056 5108 141108 5160
rect 206192 5108 206244 5160
rect 30104 5040 30156 5092
rect 127164 5040 127216 5092
rect 147680 5040 147732 5092
rect 294880 5040 294932 5092
rect 15936 4972 15988 5024
rect 108304 4972 108356 5024
rect 136916 4972 136968 5024
rect 145932 4972 145984 5024
rect 154396 4972 154448 5024
rect 364616 4972 364668 5024
rect 436836 4972 436888 5024
rect 28908 4904 28960 4956
rect 127072 4904 127124 4956
rect 138388 4904 138440 4956
rect 167184 4904 167236 4956
rect 175924 4904 175976 4956
rect 433248 4904 433300 4956
rect 479340 4904 479392 4956
rect 6460 4836 6512 4888
rect 10324 4836 10376 4888
rect 13544 4836 13596 4888
rect 125784 4836 125836 4888
rect 138296 4836 138348 4888
rect 169576 4836 169628 4888
rect 170680 4836 170732 4888
rect 480536 4836 480588 4888
rect 8760 4768 8812 4820
rect 125876 4768 125928 4820
rect 138204 4768 138256 4820
rect 162492 4768 162544 4820
rect 166632 4768 166684 4820
rect 518348 4768 518400 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 122840 4088 122892 4140
rect 123484 4088 123536 4140
rect 138848 4088 138900 4140
rect 143540 4088 143592 4140
rect 143632 4088 143684 4140
rect 147036 4156 147088 4208
rect 146944 4088 146996 4140
rect 151820 4088 151872 4140
rect 161112 4088 161164 4140
rect 182548 4088 182600 4140
rect 218704 4088 218756 4140
rect 219348 4088 219400 4140
rect 123116 4020 123168 4072
rect 131212 4020 131264 4072
rect 136824 4020 136876 4072
rect 150624 4020 150676 4072
rect 152464 4020 152516 4072
rect 163688 4020 163740 4072
rect 171876 4020 171928 4072
rect 196808 4020 196860 4072
rect 87972 3884 88024 3936
rect 122840 3884 122892 3936
rect 86868 3816 86920 3868
rect 131856 3952 131908 4004
rect 140136 3952 140188 4004
rect 164884 3952 164936 4004
rect 173164 3952 173216 4004
rect 212172 3952 212224 4004
rect 124680 3884 124732 3936
rect 134524 3884 134576 3936
rect 140780 3884 140832 3936
rect 200304 3884 200356 3936
rect 83280 3748 83332 3800
rect 123116 3748 123168 3800
rect 79692 3680 79744 3732
rect 131304 3816 131356 3868
rect 138756 3816 138808 3868
rect 140872 3816 140924 3868
rect 203892 3816 203944 3868
rect 146944 3748 146996 3800
rect 147036 3748 147088 3800
rect 232228 3748 232280 3800
rect 251180 3748 251232 3800
rect 252376 3748 252428 3800
rect 123300 3680 123352 3732
rect 130660 3680 130712 3732
rect 135168 3680 135220 3732
rect 69112 3612 69164 3664
rect 126244 3612 126296 3664
rect 127072 3612 127124 3664
rect 130292 3612 130344 3664
rect 136548 3612 136600 3664
rect 146300 3680 146352 3732
rect 267740 3680 267792 3732
rect 276020 3680 276072 3732
rect 276756 3680 276808 3732
rect 284300 3680 284352 3732
rect 285036 3680 285088 3732
rect 35900 3544 35952 3596
rect 36820 3544 36872 3596
rect 65524 3544 65576 3596
rect 123300 3544 123352 3596
rect 17040 3476 17092 3528
rect 126428 3544 126480 3596
rect 129372 3544 129424 3596
rect 130476 3544 130528 3596
rect 135444 3544 135496 3596
rect 140044 3544 140096 3596
rect 123484 3476 123536 3528
rect 124864 3476 124916 3528
rect 126980 3476 127032 3528
rect 128176 3476 128228 3528
rect 135720 3476 135772 3528
rect 138848 3476 138900 3528
rect 161296 3612 161348 3664
rect 163780 3612 163832 3664
rect 324320 3612 324372 3664
rect 140964 3544 141016 3596
rect 207388 3544 207440 3596
rect 218060 3544 218112 3596
rect 219256 3544 219308 3596
rect 219348 3544 219400 3596
rect 437940 3544 437992 3596
rect 440240 3544 440292 3596
rect 441528 3544 441580 3596
rect 448612 3544 448664 3596
rect 449808 3544 449860 3596
rect 456892 3544 456944 3596
rect 458088 3544 458140 3596
rect 474004 3544 474056 3596
rect 144736 3476 144788 3528
rect 12348 3408 12400 3460
rect 125692 3408 125744 3460
rect 131764 3408 131816 3460
rect 135904 3408 135956 3460
rect 140136 3408 140188 3460
rect 170772 3476 170824 3528
rect 173256 3476 173308 3528
rect 175464 3476 175516 3528
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 142988 3340 143040 3392
rect 147036 3340 147088 3392
rect 139032 3272 139084 3324
rect 168380 3408 168432 3460
rect 172336 3408 172388 3460
rect 462780 3476 462832 3528
rect 465080 3476 465132 3528
rect 465908 3476 465960 3528
rect 473360 3476 473412 3528
rect 474188 3476 474240 3528
rect 574744 3544 574796 3596
rect 495900 3476 495952 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 180340 3408 180392 3460
rect 475752 3408 475804 3460
rect 481640 3408 481692 3460
rect 482468 3408 482520 3460
rect 581000 3408 581052 3460
rect 147220 3340 147272 3392
rect 155408 3340 155460 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365812 3340 365864 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415492 3340 415544 3392
rect 416688 3340 416740 3392
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 137744 3204 137796 3256
rect 147128 3204 147180 3256
rect 135812 3136 135864 3188
rect 141240 3136 141292 3188
rect 144460 3136 144512 3188
rect 153016 3136 153068 3188
rect 132960 3068 133012 3120
rect 135536 3068 135588 3120
rect 136732 3068 136784 3120
rect 148324 3068 148376 3120
rect 124128 3000 124180 3052
rect 125876 3000 125928 3052
rect 135628 3000 135680 3052
rect 137652 3000 137704 3052
rect 152740 2932 152792 2984
rect 156604 2932 156656 2984
rect 349160 1504 349212 1556
rect 350448 1504 350500 1556
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 2778 580000 2834 580009
rect 2778 579935 2780 579944
rect 2832 579935 2834 579944
rect 2780 579906 2832 579912
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3252 292602 3280 293111
rect 3240 292596 3292 292602
rect 3240 292538 3292 292544
rect 3146 267200 3202 267209
rect 3146 267135 3202 267144
rect 3160 266422 3188 267135
rect 3148 266416 3200 266422
rect 3148 266358 3200 266364
rect 3238 254144 3294 254153
rect 3238 254079 3294 254088
rect 3252 253978 3280 254079
rect 3240 253972 3292 253978
rect 3240 253914 3292 253920
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3252 240174 3280 241023
rect 3240 240168 3292 240174
rect 3240 240110 3292 240116
rect 3238 228032 3294 228041
rect 3238 227967 3294 227976
rect 3252 227798 3280 227967
rect 3240 227792 3292 227798
rect 3240 227734 3292 227740
rect 3238 214976 3294 214985
rect 3238 214911 3294 214920
rect 3252 213994 3280 214911
rect 3240 213988 3292 213994
rect 3240 213930 3292 213936
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3160 187746 3188 188799
rect 3148 187740 3200 187746
rect 3148 187682 3200 187688
rect 3148 162920 3200 162926
rect 3146 162888 3148 162897
rect 3200 162888 3202 162897
rect 3146 162823 3202 162832
rect 3252 151814 3280 201855
rect 3068 151786 3280 151814
rect 3068 148374 3096 151786
rect 3344 149954 3372 306167
rect 3160 149926 3372 149954
rect 3056 148368 3108 148374
rect 3056 148310 3108 148316
rect 3160 136610 3188 149926
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 149122 3372 149767
rect 3332 149116 3384 149122
rect 3332 149058 3384 149064
rect 3240 139460 3292 139466
rect 3240 139402 3292 139408
rect 3148 136604 3200 136610
rect 3148 136546 3200 136552
rect 3148 111512 3200 111518
rect 3148 111454 3200 111460
rect 3160 110673 3188 111454
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3252 97617 3280 139402
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 3436 78985 3464 658135
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 527912 3570 527921
rect 3514 527847 3516 527856
rect 3568 527847 3570 527856
rect 3516 527818 3568 527824
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3528 474774 3556 475623
rect 3516 474768 3568 474774
rect 3516 474710 3568 474716
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3528 79626 3556 449511
rect 3516 79620 3568 79626
rect 3516 79562 3568 79568
rect 3620 79121 3648 606047
rect 3790 553888 3846 553897
rect 3790 553823 3846 553832
rect 3698 397488 3754 397497
rect 3698 397423 3754 397432
rect 3712 79762 3740 397423
rect 3700 79756 3752 79762
rect 3700 79698 3752 79704
rect 3804 79257 3832 553823
rect 3974 501800 4030 501809
rect 3974 501735 4030 501744
rect 3882 345400 3938 345409
rect 3882 345335 3938 345344
rect 3896 79898 3924 345335
rect 3884 79892 3936 79898
rect 3884 79834 3936 79840
rect 3988 79393 4016 501735
rect 4066 358456 4122 358465
rect 4066 358391 4122 358400
rect 4080 128314 4108 358391
rect 4068 128308 4120 128314
rect 4068 128250 4120 128256
rect 4816 110430 4844 683674
rect 4896 579964 4948 579970
rect 4896 579906 4948 579912
rect 4908 111790 4936 579906
rect 6184 120148 6236 120154
rect 6184 120090 6236 120096
rect 4896 111784 4948 111790
rect 4896 111726 4948 111732
rect 6196 111518 6224 120090
rect 6184 111512 6236 111518
rect 6184 111454 6236 111460
rect 4804 110424 4856 110430
rect 4804 110366 4856 110372
rect 6932 79529 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 18604 670744 18656 670750
rect 18604 670686 18656 670692
rect 7564 632120 7616 632126
rect 7564 632062 7616 632068
rect 7576 111722 7604 632062
rect 8944 527876 8996 527882
rect 8944 527818 8996 527824
rect 7656 123480 7708 123486
rect 7656 123422 7708 123428
rect 7564 111716 7616 111722
rect 7564 111658 7616 111664
rect 6918 79520 6974 79529
rect 6918 79455 6974 79464
rect 3974 79384 4030 79393
rect 3974 79319 4030 79328
rect 3790 79248 3846 79257
rect 3790 79183 3846 79192
rect 3606 79112 3662 79121
rect 3606 79047 3662 79056
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 6920 76560 6972 76566
rect 6920 76502 6972 76508
rect 2778 75304 2834 75313
rect 2778 75239 2834 75248
rect 1398 75168 1454 75177
rect 1398 75103 1454 75112
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 542 -960 654 480
rect 1412 354 1440 75103
rect 2792 16574 2820 75239
rect 4160 74044 4212 74050
rect 4160 73986 4212 73992
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 32564 3476 32570
rect 3424 32506 3476 32512
rect 3436 32473 3464 32506
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 19417 3372 24074
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3330 19408 3386 19417
rect 3330 19343 3386 19352
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 3436 6497 3464 23122
rect 4172 16574 4200 73986
rect 6932 16574 6960 76502
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4080 480 4108 4791
rect 5276 480 5304 16546
rect 6460 4888 6512 4894
rect 6460 4830 6512 4836
rect 6472 480 6500 4830
rect 7484 3482 7512 16546
rect 7576 4146 7604 36518
rect 7668 32570 7696 123422
rect 8956 113150 8984 527818
rect 13084 474768 13136 474774
rect 13084 474710 13136 474716
rect 10324 422340 10376 422346
rect 10324 422282 10376 422288
rect 10336 115938 10364 422282
rect 11704 292596 11756 292602
rect 11704 292538 11756 292544
rect 10324 115932 10376 115938
rect 10324 115874 10376 115880
rect 8944 113144 8996 113150
rect 8944 113086 8996 113092
rect 11716 80034 11744 292538
rect 13096 114510 13124 474710
rect 14464 371272 14516 371278
rect 14464 371214 14516 371220
rect 14476 117298 14504 371214
rect 17224 266416 17276 266422
rect 17224 266358 17276 266364
rect 17236 118658 17264 266358
rect 18616 135250 18644 670686
rect 21364 618316 21416 618322
rect 21364 618258 21416 618264
rect 18604 135244 18656 135250
rect 18604 135186 18656 135192
rect 21376 133890 21404 618258
rect 22744 462392 22796 462398
rect 22744 462334 22796 462340
rect 21364 133884 21416 133890
rect 21364 133826 21416 133832
rect 22756 131102 22784 462334
rect 23492 136542 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 31024 565888 31076 565894
rect 31024 565830 31076 565836
rect 28264 409896 28316 409902
rect 28264 409838 28316 409844
rect 26884 318844 26936 318850
rect 26884 318786 26936 318792
rect 25504 253972 25556 253978
rect 25504 253914 25556 253920
rect 25516 146946 25544 253914
rect 25504 146940 25556 146946
rect 25504 146882 25556 146888
rect 23480 136536 23532 136542
rect 23480 136478 23532 136484
rect 22744 131096 22796 131102
rect 22744 131038 22796 131044
rect 17316 122120 17368 122126
rect 17316 122062 17368 122068
rect 17224 118652 17276 118658
rect 17224 118594 17276 118600
rect 14464 117292 14516 117298
rect 14464 117234 14516 117240
rect 13084 114504 13136 114510
rect 13084 114446 13136 114452
rect 11704 80028 11756 80034
rect 11704 79970 11756 79976
rect 10322 77888 10378 77897
rect 10322 77823 10378 77832
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 4762
rect 9968 480 9996 8910
rect 10336 4894 10364 77823
rect 17328 71738 17356 122062
rect 26896 117230 26924 318786
rect 28276 129742 28304 409838
rect 31036 132462 31064 565830
rect 32404 514820 32456 514826
rect 32404 514762 32456 514768
rect 31024 132456 31076 132462
rect 31024 132398 31076 132404
rect 32416 132394 32444 514762
rect 32404 132388 32456 132394
rect 32404 132330 32456 132336
rect 28264 129736 28316 129742
rect 28264 129678 28316 129684
rect 26884 117224 26936 117230
rect 26884 117166 26936 117172
rect 40052 109002 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 45284 700460 45336 700466
rect 45284 700402 45336 700408
rect 44640 700392 44692 700398
rect 44640 700334 44692 700340
rect 40684 227792 40736 227798
rect 40684 227734 40736 227740
rect 40696 215966 40724 227734
rect 40684 215960 40736 215966
rect 40684 215902 40736 215908
rect 40040 108996 40092 109002
rect 40040 108938 40092 108944
rect 44652 106214 44680 700334
rect 44732 700324 44784 700330
rect 44732 700266 44784 700272
rect 44640 106208 44692 106214
rect 44640 106150 44692 106156
rect 44744 104854 44772 700266
rect 45192 261520 45244 261526
rect 45192 261462 45244 261468
rect 44916 240916 44968 240922
rect 44916 240858 44968 240864
rect 44824 240168 44876 240174
rect 44824 240110 44876 240116
rect 44732 104848 44784 104854
rect 44732 104790 44784 104796
rect 44836 78577 44864 240110
rect 44928 80481 44956 240858
rect 45008 240848 45060 240854
rect 45008 240790 45060 240796
rect 45020 141409 45048 240790
rect 45100 240780 45152 240786
rect 45100 240722 45152 240728
rect 45006 141400 45062 141409
rect 45006 141335 45062 141344
rect 45112 107642 45140 240722
rect 45204 230518 45232 261462
rect 45192 230512 45244 230518
rect 45192 230454 45244 230460
rect 45100 107636 45152 107642
rect 45100 107578 45152 107584
rect 45296 106282 45324 700402
rect 69664 396772 69716 396778
rect 69664 396714 69716 396720
rect 69676 385014 69704 396714
rect 68284 385008 68336 385014
rect 68284 384950 68336 384956
rect 69664 385008 69716 385014
rect 69664 384950 69716 384956
rect 68296 358834 68324 384950
rect 65432 358828 65484 358834
rect 65432 358770 65484 358776
rect 68284 358828 68336 358834
rect 68284 358770 68336 358776
rect 65444 358154 65472 358770
rect 64144 358148 64196 358154
rect 64144 358090 64196 358096
rect 65432 358148 65484 358154
rect 65432 358090 65484 358096
rect 45836 349852 45888 349858
rect 45836 349794 45888 349800
rect 45744 284368 45796 284374
rect 45744 284310 45796 284316
rect 45652 263628 45704 263634
rect 45652 263570 45704 263576
rect 45560 249484 45612 249490
rect 45560 249426 45612 249432
rect 45572 241514 45600 249426
rect 45480 241486 45600 241514
rect 45480 241398 45508 241486
rect 45468 241392 45520 241398
rect 45468 241334 45520 241340
rect 45468 239760 45520 239766
rect 45468 239702 45520 239708
rect 45376 238808 45428 238814
rect 45376 238750 45428 238756
rect 45388 231130 45416 238750
rect 45480 232778 45508 239702
rect 45664 232966 45692 263570
rect 45756 238814 45784 284310
rect 45848 248414 45876 349794
rect 64156 319462 64184 358090
rect 62764 319456 62816 319462
rect 62764 319398 62816 319404
rect 64144 319456 64196 319462
rect 64144 319398 64196 319404
rect 58624 315308 58676 315314
rect 58624 315250 58676 315256
rect 58636 298790 58664 315250
rect 62776 299470 62804 319398
rect 62856 305652 62908 305658
rect 62856 305594 62908 305600
rect 61476 299464 61528 299470
rect 61476 299406 61528 299412
rect 62764 299464 62816 299470
rect 62764 299406 62816 299412
rect 54484 298784 54536 298790
rect 54484 298726 54536 298732
rect 58624 298784 58676 298790
rect 58624 298726 58676 298732
rect 54496 284374 54524 298726
rect 61200 294092 61252 294098
rect 61200 294034 61252 294040
rect 60004 294024 60056 294030
rect 60004 293966 60056 293972
rect 59544 289740 59596 289746
rect 59544 289682 59596 289688
rect 59556 284374 59584 289682
rect 54484 284368 54536 284374
rect 54484 284310 54536 284316
rect 57336 284368 57388 284374
rect 57336 284310 57388 284316
rect 59544 284368 59596 284374
rect 59544 284310 59596 284316
rect 57348 280838 57376 284310
rect 60016 282946 60044 293966
rect 61212 289746 61240 294034
rect 61488 294030 61516 299406
rect 62868 294098 62896 305594
rect 68284 295384 68336 295390
rect 68284 295326 68336 295332
rect 62856 294092 62908 294098
rect 62856 294034 62908 294040
rect 61476 294024 61528 294030
rect 61476 293966 61528 293972
rect 61200 289740 61252 289746
rect 61200 289682 61252 289688
rect 68296 285734 68324 295326
rect 65708 285728 65760 285734
rect 65708 285670 65760 285676
rect 68284 285728 68336 285734
rect 68284 285670 68336 285676
rect 57980 282940 58032 282946
rect 57980 282882 58032 282888
rect 60004 282940 60056 282946
rect 60004 282882 60056 282888
rect 53104 280832 53156 280838
rect 53104 280774 53156 280780
rect 57336 280832 57388 280838
rect 57336 280774 57388 280780
rect 53116 276078 53144 280774
rect 57992 280242 58020 282882
rect 57900 280214 58020 280242
rect 57900 278798 57928 280214
rect 53840 278792 53892 278798
rect 53840 278734 53892 278740
rect 57888 278792 57940 278798
rect 57888 278734 57940 278740
rect 51724 276072 51776 276078
rect 51724 276014 51776 276020
rect 53104 276072 53156 276078
rect 53104 276014 53156 276020
rect 47584 271176 47636 271182
rect 47584 271118 47636 271124
rect 47596 263634 47624 271118
rect 47584 263628 47636 263634
rect 47584 263570 47636 263576
rect 51736 253230 51764 276014
rect 53852 271182 53880 278734
rect 65720 277438 65748 285670
rect 61384 277432 61436 277438
rect 61384 277374 61436 277380
rect 65708 277432 65760 277438
rect 65708 277374 65760 277380
rect 53840 271176 53892 271182
rect 53840 271118 53892 271124
rect 61396 261526 61424 277374
rect 61384 261520 61436 261526
rect 61384 261462 61436 261468
rect 48228 253224 48280 253230
rect 48228 253166 48280 253172
rect 51724 253224 51776 253230
rect 51724 253166 51776 253172
rect 48240 249490 48268 253166
rect 48228 249484 48280 249490
rect 48228 249426 48280 249432
rect 45848 248386 45968 248414
rect 45836 241392 45888 241398
rect 45836 241334 45888 241340
rect 45744 238808 45796 238814
rect 45744 238750 45796 238756
rect 45848 233170 45876 241334
rect 45940 239766 45968 248386
rect 71792 240922 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 86224 419552 86276 419558
rect 86224 419494 86276 419500
rect 86236 410174 86264 419494
rect 83464 410168 83516 410174
rect 83464 410110 83516 410116
rect 86224 410168 86276 410174
rect 86224 410110 86276 410116
rect 83476 371278 83504 410110
rect 77944 371272 77996 371278
rect 77944 371214 77996 371220
rect 83464 371272 83516 371278
rect 83464 371214 83516 371220
rect 77956 349858 77984 371214
rect 79324 355360 79376 355366
rect 79324 355302 79376 355308
rect 77944 349852 77996 349858
rect 77944 349794 77996 349800
rect 76564 333260 76616 333266
rect 76564 333202 76616 333208
rect 76576 321434 76604 333202
rect 79336 329594 79364 355302
rect 76656 329588 76708 329594
rect 76656 329530 76708 329536
rect 79324 329588 79376 329594
rect 79324 329530 79376 329536
rect 72424 321428 72476 321434
rect 72424 321370 72476 321376
rect 76564 321428 76616 321434
rect 76564 321370 76616 321376
rect 72436 315314 72464 321370
rect 76668 319054 76696 329530
rect 73804 319048 73856 319054
rect 73804 318990 73856 318996
rect 76656 319048 76708 319054
rect 76656 318990 76708 318996
rect 72424 315308 72476 315314
rect 72424 315250 72476 315256
rect 73816 295390 73844 318990
rect 73804 295384 73856 295390
rect 73804 295326 73856 295332
rect 71780 240916 71832 240922
rect 71780 240858 71832 240864
rect 88352 240854 88380 702406
rect 102784 502988 102836 502994
rect 102784 502930 102836 502936
rect 102796 498234 102824 502930
rect 100024 498228 100076 498234
rect 100024 498170 100076 498176
rect 102784 498228 102836 498234
rect 102784 498170 102836 498176
rect 100036 464778 100064 498170
rect 97264 464772 97316 464778
rect 97264 464714 97316 464720
rect 100024 464772 100076 464778
rect 100024 464714 100076 464720
rect 97276 458862 97304 464714
rect 88984 458856 89036 458862
rect 88984 458798 89036 458804
rect 97264 458856 97316 458862
rect 97264 458798 97316 458804
rect 88996 419558 89024 458798
rect 88984 419552 89036 419558
rect 88984 419494 89036 419500
rect 102048 384328 102100 384334
rect 102048 384270 102100 384276
rect 102060 377806 102088 384270
rect 98644 377800 98696 377806
rect 98644 377742 98696 377748
rect 102048 377800 102100 377806
rect 102048 377742 102100 377748
rect 98656 358086 98684 377742
rect 92480 358080 92532 358086
rect 92480 358022 92532 358028
rect 98644 358080 98696 358086
rect 98644 358022 98696 358028
rect 92492 355366 92520 358022
rect 92480 355360 92532 355366
rect 92480 355302 92532 355308
rect 104532 338292 104584 338298
rect 104532 338234 104584 338240
rect 104544 335374 104572 338234
rect 100760 335368 100812 335374
rect 100760 335310 100812 335316
rect 104532 335368 104584 335374
rect 104532 335310 104584 335316
rect 100772 333266 100800 335310
rect 100760 333260 100812 333266
rect 100760 333202 100812 333208
rect 88340 240848 88392 240854
rect 88340 240790 88392 240796
rect 104912 240786 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 135904 644428 135956 644434
rect 135904 644370 135956 644376
rect 135916 630698 135944 644370
rect 133144 630692 133196 630698
rect 133144 630634 133196 630640
rect 135904 630692 135956 630698
rect 135904 630634 135956 630640
rect 133156 623830 133184 630634
rect 129740 623824 129792 623830
rect 129740 623766 129792 623772
rect 133144 623824 133196 623830
rect 133144 623766 133196 623772
rect 129752 621042 129780 623766
rect 129004 621036 129056 621042
rect 129004 620978 129056 620984
rect 129740 621036 129792 621042
rect 129740 620978 129792 620984
rect 127624 598868 127676 598874
rect 127624 598810 127676 598816
rect 127636 581670 127664 598810
rect 124864 581664 124916 581670
rect 124864 581606 124916 581612
rect 127624 581664 127676 581670
rect 127624 581606 127676 581612
rect 124220 520260 124272 520266
rect 124220 520202 124272 520208
rect 122104 518968 122156 518974
rect 122104 518910 122156 518916
rect 122116 511902 122144 518910
rect 124232 514826 124260 520202
rect 124876 518974 124904 581606
rect 129016 540938 129044 620978
rect 130384 609272 130436 609278
rect 130384 609214 130436 609220
rect 130396 598874 130424 609214
rect 130384 598868 130436 598874
rect 130384 598810 130436 598816
rect 135904 550588 135956 550594
rect 135904 550530 135956 550536
rect 127624 540932 127676 540938
rect 127624 540874 127676 540880
rect 129004 540932 129056 540938
rect 129004 540874 129056 540880
rect 127636 529922 127664 540874
rect 126244 529916 126296 529922
rect 126244 529858 126296 529864
rect 127624 529916 127676 529922
rect 127624 529858 127676 529864
rect 126256 520266 126284 529858
rect 126244 520260 126296 520266
rect 126244 520202 126296 520208
rect 124864 518968 124916 518974
rect 124864 518910 124916 518916
rect 123484 514820 123536 514826
rect 123484 514762 123536 514768
rect 124220 514820 124272 514826
rect 124220 514762 124272 514768
rect 118976 511896 119028 511902
rect 118976 511838 119028 511844
rect 122104 511896 122156 511902
rect 122104 511838 122156 511844
rect 118988 507890 119016 511838
rect 116032 507884 116084 507890
rect 116032 507826 116084 507832
rect 118976 507884 119028 507890
rect 118976 507826 119028 507832
rect 116044 502994 116072 507826
rect 116032 502988 116084 502994
rect 116032 502930 116084 502936
rect 120724 453348 120776 453354
rect 120724 453290 120776 453296
rect 113824 422952 113876 422958
rect 113824 422894 113876 422900
rect 113836 384334 113864 422894
rect 119344 401668 119396 401674
rect 119344 401610 119396 401616
rect 119356 398886 119384 401610
rect 116584 398880 116636 398886
rect 116584 398822 116636 398828
rect 119344 398880 119396 398886
rect 119344 398822 119396 398828
rect 113824 384328 113876 384334
rect 113824 384270 113876 384276
rect 116596 370802 116624 398822
rect 114928 370796 114980 370802
rect 114928 370738 114980 370744
rect 116584 370796 116636 370802
rect 116584 370738 116636 370744
rect 114940 367810 114968 370738
rect 112444 367804 112496 367810
rect 112444 367746 112496 367752
rect 114928 367804 114980 367810
rect 114928 367746 114980 367752
rect 112456 353326 112484 367746
rect 120736 362982 120764 453290
rect 123496 420238 123524 514762
rect 135916 425746 135944 550530
rect 125508 425740 125560 425746
rect 125508 425682 125560 425688
rect 135904 425740 135956 425746
rect 135904 425682 135956 425688
rect 125520 422958 125548 425682
rect 125508 422952 125560 422958
rect 125508 422894 125560 422900
rect 122104 420232 122156 420238
rect 122104 420174 122156 420180
rect 123484 420232 123536 420238
rect 123484 420174 123536 420180
rect 122116 401674 122144 420174
rect 122104 401668 122156 401674
rect 122104 401610 122156 401616
rect 136652 396778 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 153212 678094 153240 702406
rect 170324 700466 170352 703520
rect 170312 700460 170364 700466
rect 170312 700402 170364 700408
rect 202800 699718 202828 703520
rect 198740 699712 198792 699718
rect 198740 699654 198792 699660
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 198752 694822 198780 699654
rect 187976 694816 188028 694822
rect 187976 694758 188028 694764
rect 198740 694816 198792 694822
rect 198740 694758 198792 694764
rect 187988 691422 188016 694758
rect 185584 691416 185636 691422
rect 185584 691358 185636 691364
rect 187976 691416 188028 691422
rect 187976 691358 188028 691364
rect 147772 678088 147824 678094
rect 147772 678030 147824 678036
rect 153200 678088 153252 678094
rect 153200 678030 153252 678036
rect 147784 675578 147812 678030
rect 147036 675572 147088 675578
rect 147036 675514 147088 675520
rect 147772 675572 147824 675578
rect 147772 675514 147824 675520
rect 147048 667894 147076 675514
rect 145564 667888 145616 667894
rect 145564 667830 145616 667836
rect 147036 667888 147088 667894
rect 147036 667830 147088 667836
rect 145576 658034 145604 667830
rect 142804 658028 142856 658034
rect 142804 657970 142856 657976
rect 145564 658028 145616 658034
rect 145564 657970 145616 657976
rect 142816 652798 142844 657970
rect 185596 653410 185624 691358
rect 177856 653404 177908 653410
rect 177856 653346 177908 653352
rect 185584 653404 185636 653410
rect 185584 653346 185636 653352
rect 142804 652792 142856 652798
rect 142804 652734 142856 652740
rect 138388 652724 138440 652730
rect 138388 652666 138440 652672
rect 138400 644502 138428 652666
rect 177868 646746 177896 653346
rect 174820 646740 174872 646746
rect 174820 646682 174872 646688
rect 177856 646740 177908 646746
rect 177856 646682 177908 646688
rect 138388 644496 138440 644502
rect 138388 644438 138440 644444
rect 174832 638246 174860 646682
rect 218072 638926 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 267660 699718 267688 703520
rect 283852 700398 283880 703520
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 293960 700392 294012 700398
rect 293960 700334 294012 700340
rect 258724 699712 258776 699718
rect 258724 699654 258776 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 258736 681834 258764 699654
rect 293972 693462 294000 700334
rect 300136 700330 300164 703520
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 396448 700392 396500 700398
rect 396448 700334 396500 700340
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 293960 693456 294012 693462
rect 293960 693398 294012 693404
rect 305644 693456 305696 693462
rect 305644 693398 305696 693404
rect 253940 681828 253992 681834
rect 253940 681770 253992 681776
rect 258724 681828 258776 681834
rect 258724 681770 258776 681776
rect 253952 678298 253980 681770
rect 305656 679658 305684 693398
rect 305644 679652 305696 679658
rect 305644 679594 305696 679600
rect 322204 679652 322256 679658
rect 322204 679594 322256 679600
rect 239404 678292 239456 678298
rect 239404 678234 239456 678240
rect 253940 678292 253992 678298
rect 253940 678234 253992 678240
rect 239416 671226 239444 678234
rect 236644 671220 236696 671226
rect 236644 671162 236696 671168
rect 239404 671220 239456 671226
rect 239404 671162 239456 671168
rect 236656 662454 236684 671162
rect 231308 662448 231360 662454
rect 231308 662390 231360 662396
rect 236644 662448 236696 662454
rect 236644 662390 236696 662396
rect 231320 659802 231348 662390
rect 224224 659796 224276 659802
rect 224224 659738 224276 659744
rect 231308 659796 231360 659802
rect 231308 659738 231360 659744
rect 214564 638920 214616 638926
rect 214564 638862 214616 638868
rect 218060 638920 218112 638926
rect 218060 638862 218112 638868
rect 152464 638240 152516 638246
rect 152464 638182 152516 638188
rect 174820 638240 174872 638246
rect 174820 638182 174872 638188
rect 152476 594862 152504 638182
rect 214576 632126 214604 638862
rect 210424 632120 210476 632126
rect 210424 632062 210476 632068
rect 214564 632120 214616 632126
rect 214564 632062 214616 632068
rect 196624 620288 196676 620294
rect 196624 620230 196676 620236
rect 196636 605130 196664 620230
rect 210436 611930 210464 632062
rect 224236 623082 224264 659738
rect 214564 623076 214616 623082
rect 214564 623018 214616 623024
rect 224224 623076 224276 623082
rect 224224 623018 224276 623024
rect 214576 620294 214604 623018
rect 322216 622470 322244 679594
rect 322204 622464 322256 622470
rect 322204 622406 322256 622412
rect 324964 622464 325016 622470
rect 324964 622406 325016 622412
rect 214564 620288 214616 620294
rect 214564 620230 214616 620236
rect 207020 611924 207072 611930
rect 207020 611866 207072 611872
rect 210424 611924 210476 611930
rect 210424 611866 210476 611872
rect 207032 609278 207060 611866
rect 207020 609272 207072 609278
rect 207020 609214 207072 609220
rect 189080 605124 189132 605130
rect 189080 605066 189132 605072
rect 196624 605124 196676 605130
rect 196624 605066 196676 605072
rect 189092 600506 189120 605066
rect 181444 600500 181496 600506
rect 181444 600442 181496 600448
rect 189080 600500 189132 600506
rect 189080 600442 189132 600448
rect 149336 594856 149388 594862
rect 149336 594798 149388 594804
rect 152464 594856 152516 594862
rect 152464 594798 152516 594804
rect 149348 592074 149376 594798
rect 146944 592068 146996 592074
rect 146944 592010 146996 592016
rect 149336 592068 149388 592074
rect 149336 592010 149388 592016
rect 146956 565146 146984 592010
rect 181456 589966 181484 600442
rect 159364 589960 159416 589966
rect 159364 589902 159416 589908
rect 181444 589960 181496 589966
rect 181444 589902 181496 589908
rect 141424 565140 141476 565146
rect 141424 565082 141476 565088
rect 146944 565140 146996 565146
rect 146944 565082 146996 565088
rect 141436 554810 141464 565082
rect 138020 554804 138072 554810
rect 138020 554746 138072 554752
rect 141424 554804 141476 554810
rect 141424 554746 141476 554752
rect 138032 550594 138060 554746
rect 138020 550588 138072 550594
rect 138020 550530 138072 550536
rect 159376 542570 159404 589902
rect 324976 570654 325004 622406
rect 324964 570648 325016 570654
rect 324964 570590 325016 570596
rect 329104 570648 329156 570654
rect 329104 570590 329156 570596
rect 155224 542564 155276 542570
rect 155224 542506 155276 542512
rect 159364 542564 159416 542570
rect 159364 542506 159416 542512
rect 155236 480350 155264 542506
rect 329116 532710 329144 570590
rect 329104 532704 329156 532710
rect 329104 532646 329156 532652
rect 331220 532704 331272 532710
rect 331220 532646 331272 532652
rect 331232 529242 331260 532646
rect 331220 529236 331272 529242
rect 331220 529178 331272 529184
rect 341524 529236 341576 529242
rect 341524 529178 341576 529184
rect 341536 517954 341564 529178
rect 341524 517948 341576 517954
rect 341524 517890 341576 517896
rect 343640 517948 343692 517954
rect 343640 517890 343692 517896
rect 343652 513330 343680 517890
rect 343640 513324 343692 513330
rect 343640 513266 343692 513272
rect 347044 513324 347096 513330
rect 347044 513266 347096 513272
rect 152464 480344 152516 480350
rect 152464 480286 152516 480292
rect 155224 480344 155276 480350
rect 155224 480286 155276 480292
rect 152476 468518 152504 480286
rect 347056 476066 347084 513266
rect 347044 476060 347096 476066
rect 347044 476002 347096 476008
rect 353300 476060 353352 476066
rect 353300 476002 353352 476008
rect 353312 472462 353340 476002
rect 353300 472456 353352 472462
rect 353300 472398 353352 472404
rect 356060 472456 356112 472462
rect 356060 472398 356112 472404
rect 142804 468512 142856 468518
rect 142804 468454 142856 468460
rect 152464 468512 152516 468518
rect 152464 468454 152516 468460
rect 142816 453354 142844 468454
rect 356072 467770 356100 472398
rect 356060 467764 356112 467770
rect 356060 467706 356112 467712
rect 359004 467764 359056 467770
rect 359004 467706 359056 467712
rect 359016 464370 359044 467706
rect 359004 464364 359056 464370
rect 359004 464306 359056 464312
rect 370504 464364 370556 464370
rect 370504 464306 370556 464312
rect 370516 459542 370544 464306
rect 370504 459536 370556 459542
rect 370504 459478 370556 459484
rect 376300 459536 376352 459542
rect 376300 459478 376352 459484
rect 376312 456414 376340 459478
rect 376300 456408 376352 456414
rect 376300 456350 376352 456356
rect 381544 456408 381596 456414
rect 381544 456350 381596 456356
rect 142804 453348 142856 453354
rect 142804 453290 142856 453296
rect 381556 437442 381584 456350
rect 381544 437436 381596 437442
rect 381544 437378 381596 437384
rect 384304 437436 384356 437442
rect 384304 437378 384356 437384
rect 384316 415410 384344 437378
rect 384304 415404 384356 415410
rect 384304 415346 384356 415352
rect 387708 415404 387760 415410
rect 387708 415346 387760 415352
rect 387720 411942 387748 415346
rect 387708 411936 387760 411942
rect 387708 411878 387760 411884
rect 136640 396772 136692 396778
rect 136640 396714 136692 396720
rect 117320 362976 117372 362982
rect 117320 362918 117372 362924
rect 120724 362976 120776 362982
rect 120724 362918 120776 362924
rect 117332 357066 117360 362918
rect 113180 357060 113232 357066
rect 113180 357002 113232 357008
rect 117320 357060 117372 357066
rect 117320 357002 117372 357008
rect 111064 353320 111116 353326
rect 111064 353262 111116 353268
rect 112444 353320 112496 353326
rect 112444 353262 112496 353268
rect 106924 348764 106976 348770
rect 106924 348706 106976 348712
rect 106936 338298 106964 348706
rect 111076 343670 111104 353262
rect 113192 348770 113220 357002
rect 113180 348764 113232 348770
rect 113180 348706 113232 348712
rect 109776 343664 109828 343670
rect 109776 343606 109828 343612
rect 111064 343664 111116 343670
rect 111064 343606 111116 343612
rect 109788 340066 109816 343606
rect 108304 340060 108356 340066
rect 108304 340002 108356 340008
rect 109776 340060 109828 340066
rect 109776 340002 109828 340008
rect 106924 338292 106976 338298
rect 106924 338234 106976 338240
rect 108316 305658 108344 340002
rect 108304 305652 108356 305658
rect 108304 305594 108356 305600
rect 104900 240780 104952 240786
rect 104900 240722 104952 240728
rect 45928 239760 45980 239766
rect 45928 239702 45980 239708
rect 45836 233164 45888 233170
rect 45836 233106 45888 233112
rect 45652 232960 45704 232966
rect 45652 232902 45704 232908
rect 73804 232960 73856 232966
rect 73804 232902 73856 232908
rect 45480 232750 45692 232778
rect 45376 231124 45428 231130
rect 45376 231066 45428 231072
rect 45664 224262 45692 232750
rect 50988 231124 51040 231130
rect 50988 231066 51040 231072
rect 46940 230512 46992 230518
rect 46940 230454 46992 230460
rect 46952 227526 46980 230454
rect 51000 228410 51028 231066
rect 50988 228404 51040 228410
rect 50988 228346 51040 228352
rect 46940 227520 46992 227526
rect 46940 227462 46992 227468
rect 50344 227520 50396 227526
rect 50344 227462 50396 227468
rect 45652 224256 45704 224262
rect 45652 224198 45704 224204
rect 48964 224256 49016 224262
rect 48964 224198 49016 224204
rect 48976 218074 49004 224198
rect 48964 218068 49016 218074
rect 48964 218010 49016 218016
rect 50356 216102 50384 227462
rect 51724 218000 51776 218006
rect 51724 217942 51776 217948
rect 50344 216096 50396 216102
rect 50344 216038 50396 216044
rect 51736 195702 51764 217942
rect 56612 195974 56640 230588
rect 58624 228404 58676 228410
rect 58624 228346 58676 228352
rect 58636 219910 58664 228346
rect 73816 224262 73844 232902
rect 116400 232416 116452 232422
rect 116400 232358 116452 232364
rect 73804 224256 73856 224262
rect 73804 224198 73856 224204
rect 77944 224256 77996 224262
rect 77944 224198 77996 224204
rect 58624 219904 58676 219910
rect 58624 219846 58676 219852
rect 64880 219904 64932 219910
rect 64880 219846 64932 219852
rect 64892 215354 64920 219846
rect 65524 216096 65576 216102
rect 65524 216038 65576 216044
rect 64880 215348 64932 215354
rect 64880 215290 64932 215296
rect 56600 195968 56652 195974
rect 56600 195910 56652 195916
rect 51724 195696 51776 195702
rect 51724 195638 51776 195644
rect 53472 195696 53524 195702
rect 53472 195638 53524 195644
rect 53484 190602 53512 195638
rect 53472 190596 53524 190602
rect 53472 190538 53524 190544
rect 55864 190596 55916 190602
rect 55864 190538 55916 190544
rect 55876 169794 55904 190538
rect 65536 177274 65564 216038
rect 68284 215348 68336 215354
rect 68284 215290 68336 215296
rect 68296 207670 68324 215290
rect 77956 215286 77984 224198
rect 77944 215280 77996 215286
rect 77944 215222 77996 215228
rect 86224 215280 86276 215286
rect 86224 215222 86276 215228
rect 68284 207664 68336 207670
rect 68284 207606 68336 207612
rect 86236 199238 86264 215222
rect 86224 199232 86276 199238
rect 86224 199174 86276 199180
rect 86972 195906 87000 230588
rect 116412 227798 116440 232358
rect 394792 232280 394844 232286
rect 394792 232222 394844 232228
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 118608 231124 118660 231130
rect 118608 231066 118660 231072
rect 116400 227792 116452 227798
rect 116400 227734 116452 227740
rect 116504 219434 116532 230588
rect 115952 219406 116532 219434
rect 90364 213988 90416 213994
rect 90364 213930 90416 213936
rect 88248 207664 88300 207670
rect 88248 207606 88300 207612
rect 88260 203590 88288 207606
rect 88248 203584 88300 203590
rect 88248 203526 88300 203532
rect 88800 199232 88852 199238
rect 88800 199174 88852 199180
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 88812 194546 88840 199174
rect 88800 194540 88852 194546
rect 88800 194482 88852 194488
rect 65524 177268 65576 177274
rect 65524 177210 65576 177216
rect 72424 177268 72476 177274
rect 72424 177210 72476 177216
rect 55864 169788 55916 169794
rect 55864 169730 55916 169736
rect 60740 169720 60792 169726
rect 60740 169662 60792 169668
rect 60752 163334 60780 169662
rect 60740 163328 60792 163334
rect 60740 163270 60792 163276
rect 66260 163328 66312 163334
rect 66260 163270 66312 163276
rect 66272 155922 66300 163270
rect 72436 156670 72464 177210
rect 86224 162920 86276 162926
rect 86224 162862 86276 162868
rect 72424 156664 72476 156670
rect 72424 156606 72476 156612
rect 79324 156664 79376 156670
rect 79324 156606 79376 156612
rect 66260 155916 66312 155922
rect 66260 155858 66312 155864
rect 67640 155916 67692 155922
rect 67640 155858 67692 155864
rect 67652 153202 67680 155858
rect 67640 153196 67692 153202
rect 67640 153138 67692 153144
rect 72424 153196 72476 153202
rect 72424 153138 72476 153144
rect 72436 141846 72464 153138
rect 79336 149734 79364 156606
rect 79324 149728 79376 149734
rect 79324 149670 79376 149676
rect 72424 141840 72476 141846
rect 72424 141782 72476 141788
rect 86236 121446 86264 162862
rect 87604 149728 87656 149734
rect 87604 149670 87656 149676
rect 86224 121440 86276 121446
rect 86224 121382 86276 121388
rect 87616 118590 87644 149670
rect 90376 126274 90404 213930
rect 112444 203584 112496 203590
rect 112444 203526 112496 203532
rect 112456 198966 112484 203526
rect 112444 198960 112496 198966
rect 112444 198902 112496 198908
rect 115204 198960 115256 198966
rect 115204 198902 115256 198908
rect 91744 194540 91796 194546
rect 91744 194482 91796 194488
rect 91756 180878 91784 194482
rect 91744 180872 91796 180878
rect 91744 180814 91796 180820
rect 95884 180872 95936 180878
rect 95884 180814 95936 180820
rect 95896 146266 95924 180814
rect 95884 146260 95936 146266
rect 95884 146202 95936 146208
rect 101404 146260 101456 146266
rect 101404 146202 101456 146208
rect 101416 137290 101444 146202
rect 101404 137284 101456 137290
rect 101404 137226 101456 137232
rect 106924 137284 106976 137290
rect 106924 137226 106976 137232
rect 90364 126268 90416 126274
rect 90364 126210 90416 126216
rect 106936 121514 106964 137226
rect 115216 130422 115244 198902
rect 115952 194614 115980 219406
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 118516 165640 118568 165646
rect 118516 165582 118568 165588
rect 118332 142860 118384 142866
rect 118332 142802 118384 142808
rect 117872 141772 117924 141778
rect 117872 141714 117924 141720
rect 116768 141024 116820 141030
rect 116768 140966 116820 140972
rect 116676 140888 116728 140894
rect 116676 140830 116728 140836
rect 116400 139596 116452 139602
rect 116400 139538 116452 139544
rect 115204 130416 115256 130422
rect 115204 130358 115256 130364
rect 116412 129742 116440 139538
rect 116584 136672 116636 136678
rect 116584 136614 116636 136620
rect 116400 129736 116452 129742
rect 116400 129678 116452 129684
rect 106924 121508 106976 121514
rect 106924 121450 106976 121456
rect 109684 121508 109736 121514
rect 109684 121450 109736 121456
rect 87604 118584 87656 118590
rect 87604 118526 87656 118532
rect 92480 118584 92532 118590
rect 92480 118526 92532 118532
rect 92492 114578 92520 118526
rect 92480 114572 92532 114578
rect 92480 114514 92532 114520
rect 95884 114572 95936 114578
rect 95884 114514 95936 114520
rect 45284 106276 45336 106282
rect 45284 106218 45336 106224
rect 95896 104786 95924 114514
rect 95884 104780 95936 104786
rect 95884 104722 95936 104728
rect 99564 104780 99616 104786
rect 99564 104722 99616 104728
rect 99576 97986 99604 104722
rect 109696 101454 109724 121450
rect 109684 101448 109736 101454
rect 109684 101390 109736 101396
rect 99564 97980 99616 97986
rect 99564 97922 99616 97928
rect 102784 97980 102836 97986
rect 102784 97922 102836 97928
rect 102796 91050 102824 97922
rect 102784 91044 102836 91050
rect 102784 90986 102836 90992
rect 105636 91044 105688 91050
rect 105636 90986 105688 90992
rect 105648 86970 105676 90986
rect 105636 86964 105688 86970
rect 105636 86906 105688 86912
rect 108120 86964 108172 86970
rect 108120 86906 108172 86912
rect 108132 80782 108160 86906
rect 108120 80776 108172 80782
rect 108120 80718 108172 80724
rect 44914 80472 44970 80481
rect 44914 80407 44970 80416
rect 116596 79150 116624 136614
rect 116688 131102 116716 140830
rect 116676 131096 116728 131102
rect 116676 131038 116728 131044
rect 116688 130121 116716 131038
rect 116674 130112 116730 130121
rect 116674 130047 116730 130056
rect 116780 128314 116808 140966
rect 117136 140956 117188 140962
rect 117136 140898 117188 140904
rect 116952 140820 117004 140826
rect 116952 140762 117004 140768
rect 116860 139528 116912 139534
rect 116860 139470 116912 139476
rect 116872 132394 116900 139470
rect 116964 132462 116992 140762
rect 117148 133890 117176 140898
rect 117780 140072 117832 140078
rect 117780 140014 117832 140020
rect 117228 139664 117280 139670
rect 117228 139606 117280 139612
rect 117240 136610 117268 139606
rect 117228 136604 117280 136610
rect 117228 136546 117280 136552
rect 117792 134722 117820 140014
rect 117884 134910 117912 141714
rect 118148 140276 118200 140282
rect 118148 140218 118200 140224
rect 117964 140208 118016 140214
rect 117964 140150 118016 140156
rect 117976 135674 118004 140150
rect 118160 135946 118188 140218
rect 118240 136536 118292 136542
rect 118240 136478 118292 136484
rect 118252 136105 118280 136478
rect 118238 136096 118294 136105
rect 118238 136031 118294 136040
rect 118160 135918 118280 135946
rect 117976 135646 118188 135674
rect 117872 134904 117924 134910
rect 117872 134846 117924 134852
rect 117792 134694 118096 134722
rect 117136 133884 117188 133890
rect 117136 133826 117188 133832
rect 117148 133498 117176 133826
rect 117148 133470 117360 133498
rect 117332 133385 117360 133470
rect 117318 133376 117374 133385
rect 117318 133311 117374 133320
rect 116952 132456 117004 132462
rect 116952 132398 117004 132404
rect 116860 132388 116912 132394
rect 116860 132330 116912 132336
rect 116872 131209 116900 132330
rect 116964 132297 116992 132398
rect 116950 132288 117006 132297
rect 116950 132223 117006 132232
rect 116858 131200 116914 131209
rect 116858 131135 116914 131144
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 129033 117360 129678
rect 117318 129024 117374 129033
rect 117318 128959 117374 128968
rect 116768 128308 116820 128314
rect 116768 128250 116820 128256
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127945 117360 128250
rect 117318 127936 117374 127945
rect 117318 127871 117374 127880
rect 117686 126848 117742 126857
rect 117686 126783 117742 126792
rect 117320 126268 117372 126274
rect 117320 126210 117372 126216
rect 117332 125769 117360 126210
rect 117318 125760 117374 125769
rect 117318 125695 117374 125704
rect 117700 122505 117728 126783
rect 117870 125760 117926 125769
rect 117870 125695 117926 125704
rect 117778 123584 117834 123593
rect 117778 123519 117834 123528
rect 117792 123486 117820 123519
rect 117780 123480 117832 123486
rect 117780 123422 117832 123428
rect 117686 122496 117742 122505
rect 117686 122431 117742 122440
rect 117700 122126 117728 122431
rect 117688 122120 117740 122126
rect 117688 122062 117740 122068
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117410 121408 117466 121417
rect 117332 120329 117360 121382
rect 117410 121343 117466 121352
rect 117318 120320 117374 120329
rect 117318 120255 117374 120264
rect 117424 120154 117452 121343
rect 117412 120148 117464 120154
rect 117412 120090 117464 120096
rect 117884 119241 117912 125695
rect 117870 119232 117926 119241
rect 117870 119167 117926 119176
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117412 117292 117464 117298
rect 117412 117234 117464 117240
rect 117320 117224 117372 117230
rect 117320 117166 117372 117172
rect 117332 117065 117360 117166
rect 117318 117056 117374 117065
rect 117318 116991 117374 117000
rect 117424 115977 117452 117234
rect 117410 115968 117466 115977
rect 117320 115932 117372 115938
rect 117410 115903 117466 115912
rect 117320 115874 117372 115880
rect 117332 114889 117360 115874
rect 117318 114880 117374 114889
rect 117318 114815 117374 114824
rect 117320 114504 117372 114510
rect 117320 114446 117372 114452
rect 117332 113801 117360 114446
rect 117318 113792 117374 113801
rect 117318 113727 117374 113736
rect 117320 113144 117372 113150
rect 117320 113086 117372 113092
rect 117332 112713 117360 113086
rect 117318 112704 117374 112713
rect 117318 112639 117374 112648
rect 117320 111784 117372 111790
rect 117320 111726 117372 111732
rect 117332 111625 117360 111726
rect 117412 111716 117464 111722
rect 117412 111658 117464 111664
rect 117318 111616 117374 111625
rect 117318 111551 117374 111560
rect 117424 110537 117452 111658
rect 117410 110528 117466 110537
rect 117410 110463 117466 110472
rect 117320 110424 117372 110430
rect 117320 110366 117372 110372
rect 117332 109449 117360 110366
rect 117318 109440 117374 109449
rect 117318 109375 117374 109384
rect 117320 108996 117372 109002
rect 117320 108938 117372 108944
rect 117332 108361 117360 108938
rect 117318 108352 117374 108361
rect 117318 108287 117374 108296
rect 117320 107636 117372 107642
rect 117320 107578 117372 107584
rect 117332 107273 117360 107578
rect 117318 107264 117374 107273
rect 117318 107199 117374 107208
rect 117320 106276 117372 106282
rect 117320 106218 117372 106224
rect 117332 106185 117360 106218
rect 117412 106208 117464 106214
rect 117318 106176 117374 106185
rect 117412 106150 117464 106156
rect 117318 106111 117374 106120
rect 117424 105097 117452 106150
rect 117410 105088 117466 105097
rect 117410 105023 117466 105032
rect 117320 104848 117372 104854
rect 117320 104790 117372 104796
rect 117332 104009 117360 104790
rect 117318 104000 117374 104009
rect 117318 103935 117374 103944
rect 118068 94217 118096 134694
rect 118054 94208 118110 94217
rect 118054 94143 118110 94152
rect 118160 92041 118188 135646
rect 118146 92032 118202 92041
rect 118146 91967 118202 91976
rect 118252 90953 118280 135918
rect 118344 93129 118372 142802
rect 118422 136640 118478 136649
rect 118422 136575 118424 136584
rect 118476 136575 118478 136584
rect 118424 136546 118476 136552
rect 118424 135244 118476 135250
rect 118424 135186 118476 135192
rect 118436 135017 118464 135186
rect 118422 135008 118478 135017
rect 118422 134943 118478 134952
rect 118424 134904 118476 134910
rect 118424 134846 118476 134852
rect 118330 93120 118386 93129
rect 118330 93055 118386 93064
rect 118238 90944 118294 90953
rect 118238 90879 118294 90888
rect 118436 89865 118464 134846
rect 118422 89856 118478 89865
rect 118422 89791 118478 89800
rect 118528 87689 118556 165582
rect 118620 102921 118648 231066
rect 146312 230574 146510 230602
rect 122104 227792 122156 227798
rect 122104 227734 122156 227740
rect 122116 214606 122144 227734
rect 122104 214600 122156 214606
rect 122104 214542 122156 214548
rect 135904 214600 135956 214606
rect 135904 214542 135956 214548
rect 118700 205692 118752 205698
rect 118700 205634 118752 205640
rect 118606 102912 118662 102921
rect 118606 102847 118662 102856
rect 118712 88777 118740 205634
rect 135916 196314 135944 214542
rect 146312 197418 146340 230574
rect 176672 229906 176700 230588
rect 174544 229900 174596 229906
rect 174544 229842 174596 229848
rect 176660 229900 176712 229906
rect 176660 229842 176712 229848
rect 166264 228472 166316 228478
rect 166264 228414 166316 228420
rect 164240 215960 164292 215966
rect 164240 215902 164292 215908
rect 154856 202156 154908 202162
rect 154856 202098 154908 202104
rect 153200 200796 153252 200802
rect 153200 200738 153252 200744
rect 148968 199436 149020 199442
rect 148968 199378 149020 199384
rect 146142 197390 146340 197418
rect 148980 197404 149008 199378
rect 153212 197470 153240 200738
rect 151084 197464 151136 197470
rect 150926 197412 151084 197418
rect 153200 197464 153252 197470
rect 150926 197406 151136 197412
rect 150926 197390 151124 197406
rect 152582 197402 152780 197418
rect 153200 197406 153252 197412
rect 154868 197402 154896 202098
rect 158904 198008 158956 198014
rect 158904 197950 158956 197956
rect 158916 197404 158944 197950
rect 152582 197396 152792 197402
rect 152582 197390 152740 197396
rect 152740 197338 152792 197344
rect 154856 197396 154908 197402
rect 154856 197338 154908 197344
rect 154488 196784 154540 196790
rect 147798 196722 147996 196738
rect 154146 196732 154488 196738
rect 154146 196726 154540 196732
rect 147798 196716 148008 196722
rect 147798 196710 147956 196716
rect 154146 196710 154528 196726
rect 147956 196658 148008 196664
rect 156144 196648 156196 196654
rect 155802 196596 156144 196602
rect 155802 196590 156196 196596
rect 155802 196574 156184 196590
rect 135904 196308 135956 196314
rect 135904 196250 135956 196256
rect 138480 196308 138532 196314
rect 138480 196250 138532 196256
rect 138112 195968 138164 195974
rect 138110 195936 138112 195945
rect 138164 195936 138166 195945
rect 138110 195871 138166 195880
rect 138492 190210 138520 196250
rect 140424 196030 140530 196058
rect 157366 196030 157564 196058
rect 140424 195945 140452 196030
rect 157536 195974 157564 196030
rect 157524 195968 157576 195974
rect 140410 195936 140466 195945
rect 139400 195900 139452 195906
rect 157524 195910 157576 195916
rect 140410 195871 140466 195880
rect 139400 195842 139452 195848
rect 139412 195537 139440 195842
rect 140778 195664 140834 195673
rect 140778 195599 140834 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 140792 194614 140820 195599
rect 140780 194608 140832 194614
rect 140780 194550 140832 194556
rect 149610 193352 149666 193361
rect 149610 193287 149666 193296
rect 140778 191856 140834 191865
rect 140778 191791 140834 191800
rect 140792 191010 140820 191791
rect 140962 191720 141018 191729
rect 140962 191655 141018 191664
rect 140870 191584 140926 191593
rect 140870 191519 140926 191528
rect 140780 191004 140832 191010
rect 140780 190946 140832 190952
rect 140778 190904 140834 190913
rect 140778 190839 140834 190848
rect 140792 190618 140820 190839
rect 140700 190590 140820 190618
rect 140700 190466 140728 190590
rect 140780 190528 140832 190534
rect 140780 190470 140832 190476
rect 140688 190460 140740 190466
rect 140688 190402 140740 190408
rect 140792 190346 140820 190470
rect 140700 190318 140820 190346
rect 138492 190182 139440 190210
rect 119344 187740 119396 187746
rect 119344 187682 119396 187688
rect 119160 141704 119212 141710
rect 119160 141646 119212 141652
rect 119068 141568 119120 141574
rect 119068 141510 119120 141516
rect 118976 141500 119028 141506
rect 118976 141442 119028 141448
rect 118884 141432 118936 141438
rect 118884 141374 118936 141380
rect 118792 140140 118844 140146
rect 118792 140082 118844 140088
rect 118804 95305 118832 140082
rect 118896 97481 118924 141374
rect 118988 98569 119016 141442
rect 119080 99657 119108 141510
rect 119172 101833 119200 141646
rect 119252 141636 119304 141642
rect 119252 141578 119304 141584
rect 119158 101824 119214 101833
rect 119158 101759 119214 101768
rect 119264 100745 119292 141578
rect 119250 100736 119306 100745
rect 119250 100671 119306 100680
rect 119066 99648 119122 99657
rect 119066 99583 119122 99592
rect 118974 98560 119030 98569
rect 118974 98495 119030 98504
rect 118882 97472 118938 97481
rect 118882 97407 118938 97416
rect 118790 95296 118846 95305
rect 118790 95231 118846 95240
rect 118698 88768 118754 88777
rect 118698 88703 118754 88712
rect 118514 87680 118570 87689
rect 118514 87615 118570 87624
rect 118514 86592 118570 86601
rect 118514 86527 118570 86536
rect 118238 84416 118294 84425
rect 118238 84351 118294 84360
rect 116584 79144 116636 79150
rect 116584 79086 116636 79092
rect 44822 78568 44878 78577
rect 44822 78503 44878 78512
rect 116584 78396 116636 78402
rect 116584 78338 116636 78344
rect 114560 78328 114612 78334
rect 114560 78270 114612 78276
rect 113824 78260 113876 78266
rect 113824 78202 113876 78208
rect 110420 78192 110472 78198
rect 110420 78134 110472 78140
rect 107660 78124 107712 78130
rect 107660 78066 107712 78072
rect 93124 78056 93176 78062
rect 93124 77998 93176 78004
rect 89720 77988 89772 77994
rect 89720 77930 89772 77936
rect 70400 76764 70452 76770
rect 70400 76706 70452 76712
rect 37278 76664 37334 76673
rect 37278 76599 37334 76608
rect 69020 76628 69072 76634
rect 20718 76528 20774 76537
rect 20718 76463 20774 76472
rect 17316 71732 17368 71738
rect 17316 71674 17368 71680
rect 13820 51740 13872 51746
rect 13820 51682 13872 51688
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11072 16574 11100 21354
rect 13832 16574 13860 51682
rect 20732 16574 20760 76463
rect 26240 75200 26292 75206
rect 26240 75142 26292 75148
rect 11072 16546 11192 16574
rect 13832 16546 14320 16574
rect 20732 16546 21864 16574
rect 10324 4888 10376 4894
rect 10324 4830 10376 4836
rect 11164 480 11192 16546
rect 13544 4888 13596 4894
rect 13544 4830 13596 4836
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12360 480 12388 3402
rect 13556 480 13584 4830
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 480 15976 4966
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 480 17080 3470
rect 18248 480 18276 6122
rect 19444 480 19472 6190
rect 20626 3360 20682 3369
rect 20626 3295 20682 3304
rect 20640 480 20668 3295
rect 21836 480 21864 16546
rect 25320 10396 25372 10402
rect 25320 10338 25372 10344
rect 24216 7608 24268 7614
rect 23018 7576 23074 7585
rect 24216 7550 24268 7556
rect 23018 7511 23074 7520
rect 23032 480 23060 7511
rect 24228 480 24256 7550
rect 25332 480 25360 10338
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 75142
rect 35898 73808 35954 73817
rect 35898 73743 35954 73752
rect 30380 44940 30432 44946
rect 30380 44882 30432 44888
rect 27620 44872 27672 44878
rect 27620 44814 27672 44820
rect 27632 16574 27660 44814
rect 30392 16574 30420 44882
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31772 16574 31800 32370
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27724 480 27752 16546
rect 30104 5092 30156 5098
rect 30104 5034 30156 5040
rect 28908 4956 28960 4962
rect 28908 4898 28960 4904
rect 28920 480 28948 4898
rect 30116 480 30144 5034
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 34796 7676 34848 7682
rect 34796 7618 34848 7624
rect 33600 6316 33652 6322
rect 33600 6258 33652 6264
rect 33612 480 33640 6258
rect 34808 480 34836 7618
rect 35912 3602 35940 73743
rect 37292 16574 37320 76599
rect 69020 76570 69072 76576
rect 51080 75404 51132 75410
rect 51080 75346 51132 75352
rect 49700 75336 49752 75342
rect 49700 75278 49752 75284
rect 46940 75268 46992 75274
rect 46940 75210 46992 75216
rect 45560 37936 45612 37942
rect 45560 37878 45612 37884
rect 38660 35216 38712 35222
rect 38660 35158 38712 35164
rect 38672 16574 38700 35158
rect 42800 18624 42852 18630
rect 42800 18566 42852 18572
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 35992 10328 36044 10334
rect 35992 10270 36044 10276
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 36004 480 36032 10270
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36832 354 36860 3538
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41878 8936 41934 8945
rect 41878 8871 41934 8880
rect 40682 6216 40738 6225
rect 40682 6151 40738 6160
rect 40696 480 40724 6151
rect 41892 480 41920 8871
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 18566
rect 45572 16574 45600 37878
rect 46952 16574 46980 75210
rect 49712 16574 49740 75278
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 45468 9036 45520 9042
rect 45468 8978 45520 8984
rect 44272 6384 44324 6390
rect 44272 6326 44324 6332
rect 44284 480 44312 6326
rect 45480 480 45508 8978
rect 46676 480 46704 16546
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 7744 49016 7750
rect 48964 7686 49016 7692
rect 48976 480 49004 7686
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 75346
rect 57978 74080 58034 74089
rect 57978 74015 58034 74024
rect 53838 73944 53894 73953
rect 53838 73879 53894 73888
rect 53852 16574 53880 73879
rect 57992 16574 58020 74015
rect 60740 73908 60792 73914
rect 60740 73850 60792 73856
rect 60752 16574 60780 73850
rect 67640 45008 67692 45014
rect 67640 44950 67692 44956
rect 63500 18692 63552 18698
rect 63500 18634 63552 18640
rect 63512 16574 63540 18634
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 60752 16546 61608 16574
rect 63512 16546 64368 16574
rect 52552 9172 52604 9178
rect 52552 9114 52604 9120
rect 52564 480 52592 9114
rect 53748 9104 53800 9110
rect 53748 9046 53800 9052
rect 53760 480 53788 9046
rect 54956 480 54984 16546
rect 57242 9208 57298 9217
rect 57242 9143 57298 9152
rect 56046 9072 56102 9081
rect 56046 9007 56102 9016
rect 56060 480 56088 9007
rect 57256 480 57284 9143
rect 58452 480 58480 16546
rect 60832 9308 60884 9314
rect 60832 9250 60884 9256
rect 59636 9240 59688 9246
rect 59636 9182 59688 9188
rect 59648 480 59676 9182
rect 60844 480 60872 9250
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63224 5160 63276 5166
rect 63224 5102 63276 5108
rect 63236 480 63264 5102
rect 64340 480 64368 16546
rect 66720 6452 66772 6458
rect 66720 6394 66772 6400
rect 65524 3596 65576 3602
rect 65524 3538 65576 3544
rect 65536 480 65564 3538
rect 66732 480 66760 6394
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 44950
rect 69032 16574 69060 76570
rect 70412 16574 70440 76706
rect 75920 75472 75972 75478
rect 75920 75414 75972 75420
rect 71778 74216 71834 74225
rect 71778 74151 71834 74160
rect 71792 16574 71820 74151
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 69112 3664 69164 3670
rect 69112 3606 69164 3612
rect 69124 480 69152 3606
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 74998 10296 75054 10305
rect 74998 10231 75054 10240
rect 73802 6352 73858 6361
rect 73802 6287 73858 6296
rect 73816 480 73844 6287
rect 75012 480 75040 10231
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 75414
rect 88340 55888 88392 55894
rect 88340 55830 88392 55836
rect 88352 16574 88380 55830
rect 89732 16574 89760 77930
rect 91098 44840 91154 44849
rect 91098 44775 91154 44784
rect 91112 16574 91140 44775
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85672 10600 85724 10606
rect 85672 10542 85724 10548
rect 81624 10532 81676 10538
rect 81624 10474 81676 10480
rect 78128 10464 78180 10470
rect 78128 10406 78180 10412
rect 77392 6520 77444 6526
rect 77392 6462 77444 6468
rect 77404 480 77432 6462
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10406
rect 80888 6588 80940 6594
rect 80888 6530 80940 6536
rect 79692 3732 79744 3738
rect 79692 3674 79744 3680
rect 79704 480 79732 3674
rect 80900 480 80928 6530
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 10474
rect 84476 7812 84528 7818
rect 84476 7754 84528 7760
rect 83280 3800 83332 3806
rect 83280 3742 83332 3748
rect 83292 480 83320 3742
rect 84488 480 84516 7754
rect 85684 480 85712 10542
rect 87972 3936 88024 3942
rect 87972 3878 88024 3884
rect 86868 3868 86920 3874
rect 86868 3810 86920 3816
rect 86880 480 86908 3810
rect 87984 480 88012 3878
rect 89180 480 89208 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92478 10432 92534 10441
rect 93136 10402 93164 77998
rect 102140 76832 102192 76838
rect 102140 76774 102192 76780
rect 93860 76696 93912 76702
rect 93860 76638 93912 76644
rect 93872 16574 93900 76638
rect 96620 72480 96672 72486
rect 96620 72422 96672 72428
rect 95240 57248 95292 57254
rect 95240 57190 95292 57196
rect 95252 16574 95280 57190
rect 96632 16574 96660 72422
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 92478 10367 92534 10376
rect 93124 10396 93176 10402
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10367
rect 93124 10338 93176 10344
rect 93952 5228 94004 5234
rect 93952 5170 94004 5176
rect 93964 480 93992 5170
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 99840 10396 99892 10402
rect 99840 10338 99892 10344
rect 98644 7880 98696 7886
rect 98644 7822 98696 7828
rect 98656 480 98684 7822
rect 99852 480 99880 10338
rect 102152 6914 102180 76774
rect 102232 61396 102284 61402
rect 102232 61338 102284 61344
rect 102244 16574 102272 61338
rect 107672 16574 107700 78066
rect 102244 16546 103376 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 101036 5296 101088 5302
rect 101036 5238 101088 5244
rect 101048 480 101076 5238
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 106464 11756 106516 11762
rect 106464 11698 106516 11704
rect 105728 7948 105780 7954
rect 105728 7890 105780 7896
rect 104532 6656 104584 6662
rect 104532 6598 104584 6604
rect 104544 480 104572 6598
rect 105740 480 105768 7890
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 11698
rect 108132 480 108160 16546
rect 109314 7712 109370 7721
rect 109314 7647 109370 7656
rect 108304 5364 108356 5370
rect 108304 5306 108356 5312
rect 108316 5030 108344 5306
rect 108304 5024 108356 5030
rect 108304 4966 108356 4972
rect 109328 480 109356 7647
rect 110432 3398 110460 78134
rect 111798 76800 111854 76809
rect 111798 76735 111854 76744
rect 111812 16574 111840 76735
rect 111812 16546 112392 16574
rect 110510 10568 110566 10577
rect 110510 10503 110566 10512
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 10503
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113836 5370 113864 78202
rect 114572 16574 114600 78270
rect 116596 37942 116624 78338
rect 118252 46918 118280 84351
rect 118330 83328 118386 83337
rect 118330 83263 118386 83272
rect 118240 46912 118292 46918
rect 118240 46854 118292 46860
rect 116584 37936 116636 37942
rect 116584 37878 116636 37884
rect 118344 22778 118372 83263
rect 118528 80646 118556 86527
rect 118606 85504 118662 85513
rect 118606 85439 118662 85448
rect 118516 80640 118568 80646
rect 118516 80582 118568 80588
rect 118620 80578 118648 85439
rect 118608 80572 118660 80578
rect 118608 80514 118660 80520
rect 119356 78033 119384 187682
rect 139412 187649 139440 190182
rect 139398 187640 139454 187649
rect 139398 187575 139454 187584
rect 140700 186130 140728 190318
rect 140780 190256 140832 190262
rect 140780 190198 140832 190204
rect 140792 186289 140820 190198
rect 140778 186280 140834 186289
rect 140778 186215 140834 186224
rect 140700 186102 140820 186130
rect 140792 182617 140820 186102
rect 140778 182608 140834 182617
rect 140778 182543 140834 182552
rect 140884 182481 140912 191519
rect 140976 182753 141004 191655
rect 149624 190534 149652 193287
rect 144736 190528 144788 190534
rect 144394 190476 144736 190482
rect 144394 190470 144788 190476
rect 149612 190528 149664 190534
rect 149612 190470 149664 190476
rect 144394 190454 144776 190470
rect 164252 189652 164280 215902
rect 166276 196790 166304 228414
rect 166264 196784 166316 196790
rect 166264 196726 166316 196732
rect 174556 196722 174584 229842
rect 180064 228404 180116 228410
rect 180064 228346 180116 228352
rect 174544 196716 174596 196722
rect 174544 196658 174596 196664
rect 165434 193352 165490 193361
rect 165434 193287 165490 193296
rect 165448 190398 165476 193287
rect 165436 190392 165488 190398
rect 165436 190334 165488 190340
rect 165436 189100 165488 189106
rect 165436 189042 165488 189048
rect 140962 182744 141018 182753
rect 140962 182679 141018 182688
rect 140870 182472 140926 182481
rect 140870 182407 140926 182416
rect 136376 182158 136758 182186
rect 136376 180130 136404 182158
rect 144460 181008 144512 181014
rect 136468 180934 136758 180962
rect 146024 181008 146076 181014
rect 144642 180976 144698 180985
rect 144460 180950 144512 180956
rect 144472 180948 144500 180950
rect 144578 180934 144642 180962
rect 121460 180124 121512 180130
rect 121460 180066 121512 180072
rect 136364 180124 136416 180130
rect 136364 180066 136416 180072
rect 121472 139890 121500 180066
rect 135996 178900 136048 178906
rect 135996 178842 136048 178848
rect 122840 178696 122892 178702
rect 122840 178638 122892 178644
rect 122852 151814 122880 178638
rect 136008 177342 136036 178842
rect 136468 178702 136496 180934
rect 144642 180911 144698 180920
rect 146022 180976 146024 180985
rect 146076 180976 146078 180985
rect 146022 180911 146078 180920
rect 136560 179982 136758 180010
rect 136560 178906 136588 179982
rect 136548 178900 136600 178906
rect 136548 178842 136600 178848
rect 136744 178786 136772 179044
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136560 178758 136772 178786
rect 141606 178800 141662 178809
rect 136456 178696 136508 178702
rect 136456 178638 136508 178644
rect 136560 178514 136588 178758
rect 141606 178735 141662 178744
rect 136192 178486 136588 178514
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 135996 177336 136048 177342
rect 135996 177278 136048 177284
rect 124232 151814 124260 177278
rect 126980 176112 127032 176118
rect 126980 176054 127032 176060
rect 125600 175976 125652 175982
rect 125600 175918 125652 175924
rect 125612 151814 125640 175918
rect 126992 151814 127020 176054
rect 136192 175982 136220 178486
rect 136284 177942 136758 177970
rect 136284 176118 136312 177942
rect 136376 176990 136758 177018
rect 136272 176112 136324 176118
rect 136272 176054 136324 176060
rect 136180 175976 136232 175982
rect 136180 175918 136232 175924
rect 136376 175234 136404 176990
rect 141620 175982 141648 178735
rect 142066 178664 142122 178673
rect 142066 178599 142122 178608
rect 141698 178528 141754 178537
rect 141698 178463 141754 178472
rect 141608 175976 141660 175982
rect 136560 175902 136758 175930
rect 141608 175918 141660 175924
rect 128360 175228 128412 175234
rect 128360 175170 128412 175176
rect 136364 175228 136416 175234
rect 136364 175170 136416 175176
rect 128372 151814 128400 175170
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 136560 173894 136588 175902
rect 131120 172576 131172 172582
rect 131120 172518 131172 172524
rect 122852 151786 122972 151814
rect 124232 151786 124536 151814
rect 125612 151786 126100 151814
rect 126992 151786 127664 151814
rect 128372 151786 129228 151814
rect 122944 139890 122972 151786
rect 124508 139890 124536 151786
rect 126072 139890 126100 151786
rect 127636 139890 127664 151786
rect 129200 139890 129228 151786
rect 131132 139890 131160 172518
rect 132500 171148 132552 171154
rect 132500 171090 132552 171096
rect 132512 139890 132540 171090
rect 133892 139890 133920 173878
rect 136560 173866 136680 173894
rect 136652 172582 136680 173866
rect 136640 172576 136692 172582
rect 136640 172518 136692 172524
rect 135260 171692 135312 171698
rect 135260 171634 135312 171640
rect 135272 151814 135300 171634
rect 136744 171154 136772 174964
rect 141712 174758 141740 178463
rect 142080 174826 142108 178599
rect 142068 174820 142120 174826
rect 142068 174762 142120 174768
rect 144104 174758 144132 178871
rect 149336 176044 149388 176050
rect 149336 175986 149388 175992
rect 144460 175568 144512 175574
rect 144460 175510 144512 175516
rect 141700 174752 141752 174758
rect 141700 174694 141752 174700
rect 144092 174752 144144 174758
rect 144092 174694 144144 174700
rect 137376 173936 137428 173942
rect 137428 173884 137586 173890
rect 137376 173878 137586 173884
rect 137388 173862 137586 173878
rect 138020 172168 138072 172174
rect 138020 172110 138072 172116
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 138032 151814 138060 172110
rect 138676 171698 138704 173196
rect 139596 173182 139702 173210
rect 138664 171692 138716 171698
rect 138664 171634 138716 171640
rect 135272 151786 135484 151814
rect 138032 151786 138612 151814
rect 135456 139890 135484 151786
rect 137744 143472 137796 143478
rect 137744 143414 137796 143420
rect 137756 139890 137784 143414
rect 121472 139862 121808 139890
rect 122944 139862 123372 139890
rect 124508 139862 124936 139890
rect 126072 139862 126500 139890
rect 127636 139862 128064 139890
rect 129200 139862 129628 139890
rect 131132 139862 131192 139890
rect 132512 139862 132756 139890
rect 133892 139862 134320 139890
rect 135456 139862 135884 139890
rect 137448 139862 137784 139890
rect 138584 139890 138612 151786
rect 139596 143478 139624 173182
rect 140792 172174 140820 173196
rect 140780 172168 140832 172174
rect 140780 172110 140832 172116
rect 139584 143472 139636 143478
rect 139584 143414 139636 143420
rect 142068 142248 142120 142254
rect 142068 142190 142120 142196
rect 140688 142180 140740 142186
rect 140688 142122 140740 142128
rect 140700 139890 140728 142122
rect 138584 139862 139012 139890
rect 140576 139862 140728 139890
rect 142080 139890 142108 142190
rect 142264 142186 142292 173196
rect 142526 172952 142582 172961
rect 142526 172887 142582 172896
rect 142436 166320 142488 166326
rect 142436 166262 142488 166268
rect 142448 142254 142476 166262
rect 142540 142934 142568 172887
rect 142632 166326 142660 173196
rect 142620 166320 142672 166326
rect 142620 166262 142672 166268
rect 143644 161474 143672 173196
rect 143552 161446 143672 161474
rect 142528 142928 142580 142934
rect 142528 142870 142580 142876
rect 142436 142248 142488 142254
rect 142436 142190 142488 142196
rect 142252 142180 142304 142186
rect 142252 142122 142304 142128
rect 143552 139890 143580 161446
rect 144472 143070 144500 175510
rect 149348 175409 149376 175986
rect 162492 175976 162544 175982
rect 162492 175918 162544 175924
rect 149980 175568 150032 175574
rect 149980 175510 150032 175516
rect 149992 175508 150020 175510
rect 154396 175432 154448 175438
rect 149334 175400 149390 175409
rect 149334 175335 149390 175344
rect 154394 175400 154396 175409
rect 154448 175400 154450 175409
rect 154394 175335 154450 175344
rect 145472 174752 145524 174758
rect 145472 174694 145524 174700
rect 144460 143064 144512 143070
rect 144460 143006 144512 143012
rect 144932 139890 144960 173196
rect 145484 143002 145512 174694
rect 152464 174684 152516 174690
rect 152464 174626 152516 174632
rect 156512 174684 156564 174690
rect 156512 174626 156564 174632
rect 152476 174570 152504 174626
rect 152398 174542 152504 174570
rect 146312 151814 146340 173196
rect 146484 166320 146536 166326
rect 146484 166262 146536 166268
rect 146312 151786 146432 151814
rect 145472 142996 145524 143002
rect 145472 142938 145524 142944
rect 146404 139890 146432 151786
rect 146496 143478 146524 166262
rect 146680 161474 146708 173196
rect 147600 166326 147628 173196
rect 149348 172990 149376 173196
rect 149336 172984 149388 172990
rect 149336 172926 149388 172932
rect 147588 166320 147640 166326
rect 147588 166262 147640 166268
rect 149624 161474 149652 173196
rect 150636 161474 150664 173196
rect 151452 172984 151504 172990
rect 151452 172926 151504 172932
rect 146588 161446 146708 161474
rect 149532 161446 149652 161474
rect 150544 161446 150664 161474
rect 146588 143546 146616 161446
rect 146576 143540 146628 143546
rect 146576 143482 146628 143488
rect 148048 143540 148100 143546
rect 148048 143482 148100 143488
rect 146484 143472 146536 143478
rect 146484 143414 146536 143420
rect 148060 139890 148088 143482
rect 149532 142186 149560 161446
rect 149612 143472 149664 143478
rect 149612 143414 149664 143420
rect 149520 142180 149572 142186
rect 149520 142122 149572 142128
rect 149624 139890 149652 143414
rect 150544 143138 150572 161446
rect 150532 143132 150584 143138
rect 150532 143074 150584 143080
rect 151464 139890 151492 172926
rect 152660 161474 152688 173196
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 152476 143478 152504 161446
rect 152464 143472 152516 143478
rect 152464 143414 152516 143420
rect 153488 143410 153516 173182
rect 155222 156632 155278 156641
rect 155222 156567 155278 156576
rect 155236 143546 155264 156567
rect 155224 143540 155276 143546
rect 155224 143482 155276 143488
rect 153476 143404 153528 143410
rect 153476 143346 153528 143352
rect 154580 143132 154632 143138
rect 154580 143074 154632 143080
rect 152740 142180 152792 142186
rect 152740 142122 152792 142128
rect 152752 139890 152780 142122
rect 154592 139890 154620 143074
rect 156524 139890 156552 174626
rect 161480 174548 161532 174554
rect 161480 174490 161532 174496
rect 159652 172990 159680 173196
rect 158444 172984 158496 172990
rect 158444 172926 158496 172932
rect 159640 172984 159692 172990
rect 159640 172926 159692 172932
rect 158456 148442 158484 172926
rect 161492 151814 161520 174490
rect 162504 172990 162532 175918
rect 165448 175545 165476 189042
rect 165434 175536 165490 175545
rect 165434 175471 165490 175480
rect 162492 172984 162544 172990
rect 162492 172926 162544 172932
rect 161492 151786 162072 151814
rect 158444 148436 158496 148442
rect 158444 148378 158496 148384
rect 160100 143540 160152 143546
rect 160100 143482 160152 143488
rect 157432 143472 157484 143478
rect 157432 143414 157484 143420
rect 142080 139862 142140 139890
rect 143552 139862 143704 139890
rect 144932 139862 145268 139890
rect 146404 139862 146832 139890
rect 148060 139862 148396 139890
rect 149624 139862 149960 139890
rect 151464 139862 151524 139890
rect 152752 139862 153088 139890
rect 154592 139862 154652 139890
rect 156216 139862 156552 139890
rect 157444 139890 157472 143414
rect 158996 143404 159048 143410
rect 158996 143346 159048 143352
rect 159008 139890 159036 143346
rect 160112 140350 160140 143482
rect 160560 143064 160612 143070
rect 160560 143006 160612 143012
rect 160100 140344 160152 140350
rect 160100 140286 160152 140292
rect 160572 139890 160600 143006
rect 162044 139890 162072 151786
rect 163516 143070 163544 175100
rect 171138 174584 171194 174593
rect 171138 174519 171194 174528
rect 167000 174344 167052 174350
rect 167000 174286 167052 174292
rect 163608 143138 163636 173196
rect 164528 173182 164634 173210
rect 163596 143132 163648 143138
rect 163596 143074 163648 143080
rect 164528 143070 164556 173182
rect 165528 172984 165580 172990
rect 165434 172952 165490 172961
rect 165528 172926 165580 172932
rect 165434 172887 165490 172896
rect 164976 148436 165028 148442
rect 164976 148378 165028 148384
rect 164988 143478 165016 148378
rect 165448 143546 165476 172887
rect 165436 143540 165488 143546
rect 165436 143482 165488 143488
rect 164976 143472 165028 143478
rect 164976 143414 165028 143420
rect 163504 143064 163556 143070
rect 163504 143006 163556 143012
rect 164516 143064 164568 143070
rect 164516 143006 164568 143012
rect 163688 142996 163740 143002
rect 163688 142938 163740 142944
rect 163700 139890 163728 142938
rect 165540 139890 165568 172926
rect 167012 139890 167040 174286
rect 171152 151814 171180 174519
rect 171152 151786 171456 151814
rect 169944 143540 169996 143546
rect 169944 143482 169996 143488
rect 168380 143472 168432 143478
rect 168380 143414 168432 143420
rect 168392 139890 168420 143414
rect 169956 139890 169984 143482
rect 171428 139890 171456 151786
rect 179420 149116 179472 149122
rect 179420 149058 179472 149064
rect 174636 143132 174688 143138
rect 174636 143074 174688 143080
rect 173072 142928 173124 142934
rect 173072 142870 173124 142876
rect 173084 139890 173112 142870
rect 174648 139890 174676 143074
rect 176200 143064 176252 143070
rect 176200 143006 176252 143012
rect 176212 139890 176240 143006
rect 178040 142996 178092 143002
rect 178040 142938 178092 142944
rect 178052 139890 178080 142938
rect 157444 139862 157780 139890
rect 159008 139862 159344 139890
rect 160572 139862 160908 139890
rect 162044 139862 162472 139890
rect 163700 139862 164036 139890
rect 165540 139862 165600 139890
rect 167012 139862 167164 139890
rect 168392 139862 168728 139890
rect 169956 139862 170292 139890
rect 171428 139862 171856 139890
rect 173084 139862 173420 139890
rect 174648 139862 174984 139890
rect 176212 139862 176548 139890
rect 178052 139862 178112 139890
rect 120540 139800 120592 139806
rect 120540 139742 120592 139748
rect 120552 135017 120580 139742
rect 120632 139732 120684 139738
rect 120632 139674 120684 139680
rect 120644 136105 120672 139674
rect 120630 136096 120686 136105
rect 120630 136031 120686 136040
rect 120538 135008 120594 135017
rect 120538 134943 120594 134952
rect 120724 130416 120776 130422
rect 120724 130358 120776 130364
rect 119436 101448 119488 101454
rect 119436 101390 119488 101396
rect 119342 78024 119398 78033
rect 119342 77959 119398 77968
rect 119448 77246 119476 101390
rect 120632 84244 120684 84250
rect 120632 84186 120684 84192
rect 120080 80776 120132 80782
rect 120080 80718 120132 80724
rect 120092 77858 120120 80718
rect 120644 79286 120672 84186
rect 120632 79280 120684 79286
rect 120632 79222 120684 79228
rect 120080 77852 120132 77858
rect 120080 77794 120132 77800
rect 119436 77240 119488 77246
rect 119436 77182 119488 77188
rect 118700 76900 118752 76906
rect 118700 76842 118752 76848
rect 118332 22772 118384 22778
rect 118332 22714 118384 22720
rect 114572 16546 114784 16574
rect 113824 5364 113876 5370
rect 113824 5306 113876 5312
rect 114008 5364 114060 5370
rect 114008 5306 114060 5312
rect 114020 480 114048 5306
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 117320 11824 117372 11830
rect 117320 11766 117372 11772
rect 116400 8016 116452 8022
rect 116400 7958 116452 7964
rect 116412 480 116440 7958
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 11766
rect 118712 3398 118740 76842
rect 120736 75954 120764 130358
rect 179432 126857 179460 149058
rect 179512 141840 179564 141846
rect 179512 141782 179564 141788
rect 179524 139874 179552 141782
rect 179512 139868 179564 139874
rect 179512 139810 179564 139816
rect 179512 139460 179564 139466
rect 179512 139402 179564 139408
rect 179524 128217 179552 139402
rect 179510 128208 179566 128217
rect 179510 128143 179566 128152
rect 179418 126848 179474 126857
rect 179418 126783 179474 126792
rect 179972 85604 180024 85610
rect 179972 85546 180024 85552
rect 178960 81252 179012 81258
rect 178960 81194 179012 81200
rect 178972 80782 179000 81194
rect 178960 80776 179012 80782
rect 178960 80718 179012 80724
rect 179984 80714 180012 85546
rect 178592 80708 178644 80714
rect 178592 80650 178644 80656
rect 179972 80708 180024 80714
rect 179972 80650 180024 80656
rect 174452 80572 174504 80578
rect 174452 80514 174504 80520
rect 174464 80442 174492 80514
rect 174452 80436 174504 80442
rect 174452 80378 174504 80384
rect 175280 80436 175332 80442
rect 175280 80378 175332 80384
rect 174452 80300 174504 80306
rect 174452 80242 174504 80248
rect 125230 80200 125286 80209
rect 174464 80170 174492 80242
rect 125230 80135 125286 80144
rect 174452 80164 174504 80170
rect 124770 79928 124826 79937
rect 123668 79892 123720 79898
rect 124770 79863 124826 79872
rect 123668 79834 123720 79840
rect 122196 78464 122248 78470
rect 122196 78406 122248 78412
rect 122102 78160 122158 78169
rect 122102 78095 122158 78104
rect 120816 77376 120868 77382
rect 120816 77318 120868 77324
rect 120724 75948 120776 75954
rect 120724 75890 120776 75896
rect 118792 73976 118844 73982
rect 118792 73918 118844 73924
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 73918
rect 120080 60240 120132 60246
rect 120080 60182 120132 60188
rect 120092 16574 120120 60182
rect 120828 32434 120856 77318
rect 121460 75540 121512 75546
rect 121460 75482 121512 75488
rect 120816 32428 120868 32434
rect 120816 32370 120868 32376
rect 120092 16546 120672 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 121472 6914 121500 75482
rect 122116 7614 122144 78095
rect 122208 35222 122236 78406
rect 122932 78192 122984 78198
rect 122932 78134 122984 78140
rect 123300 78192 123352 78198
rect 123300 78134 123352 78140
rect 122944 77518 122972 78134
rect 123312 77994 123340 78134
rect 123392 78124 123444 78130
rect 123392 78066 123444 78072
rect 123300 77988 123352 77994
rect 123300 77930 123352 77936
rect 123404 77586 123432 78066
rect 123392 77580 123444 77586
rect 123392 77522 123444 77528
rect 122932 77512 122984 77518
rect 122932 77454 122984 77460
rect 123576 77444 123628 77450
rect 123576 77386 123628 77392
rect 123484 77036 123536 77042
rect 123484 76978 123536 76984
rect 122196 35216 122248 35222
rect 122196 35158 122248 35164
rect 122104 7608 122156 7614
rect 122104 7550 122156 7556
rect 121472 6886 122328 6914
rect 122300 480 122328 6886
rect 123496 4146 123524 76978
rect 123588 60246 123616 77386
rect 123680 75313 123708 79834
rect 124036 77852 124088 77858
rect 124036 77794 124088 77800
rect 124128 77852 124180 77858
rect 124128 77794 124180 77800
rect 124048 76022 124076 77794
rect 124036 76016 124088 76022
rect 124036 75958 124088 75964
rect 123666 75304 123722 75313
rect 123666 75239 123722 75248
rect 123576 60240 123628 60246
rect 123576 60182 123628 60188
rect 122840 4140 122892 4146
rect 122840 4082 122892 4088
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 122852 3942 122880 4082
rect 123116 4072 123168 4078
rect 123116 4014 123168 4020
rect 122840 3936 122892 3942
rect 122840 3878 122892 3884
rect 123128 3806 123156 4014
rect 123116 3800 123168 3806
rect 123116 3742 123168 3748
rect 123300 3732 123352 3738
rect 123300 3674 123352 3680
rect 123312 3602 123340 3674
rect 123300 3596 123352 3602
rect 123300 3538 123352 3544
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 123496 480 123524 3470
rect 124140 3058 124168 77794
rect 124784 76566 124812 79863
rect 125048 79824 125100 79830
rect 125048 79766 125100 79772
rect 124956 77988 125008 77994
rect 124956 77930 125008 77936
rect 124864 76968 124916 76974
rect 124864 76910 124916 76916
rect 124772 76560 124824 76566
rect 124772 76502 124824 76508
rect 124772 72412 124824 72418
rect 124772 72354 124824 72360
rect 124784 70394 124812 72354
rect 124232 70366 124812 70394
rect 124232 36582 124260 70366
rect 124220 36576 124272 36582
rect 124220 36518 124272 36524
rect 124680 3936 124732 3942
rect 124680 3878 124732 3884
rect 124128 3052 124180 3058
rect 124128 2994 124180 3000
rect 124692 480 124720 3878
rect 124876 3534 124904 76910
rect 124968 6254 124996 77930
rect 125060 77897 125088 79766
rect 125140 79688 125192 79694
rect 125140 79630 125192 79636
rect 125046 77888 125102 77897
rect 125046 77823 125102 77832
rect 125152 77738 125180 79630
rect 125060 77710 125180 77738
rect 125060 55894 125088 77710
rect 125140 77648 125192 77654
rect 125140 77590 125192 77596
rect 125048 55888 125100 55894
rect 125048 55830 125100 55836
rect 125152 51746 125180 77590
rect 125244 57254 125272 80135
rect 174452 80106 174504 80112
rect 174544 80096 174596 80102
rect 125428 80022 125580 80050
rect 125322 79792 125378 79801
rect 125322 79727 125378 79736
rect 125336 78266 125364 79727
rect 125324 78260 125376 78266
rect 125324 78202 125376 78208
rect 125324 77920 125376 77926
rect 125324 77862 125376 77868
rect 125336 61402 125364 77862
rect 125428 72418 125456 80022
rect 125508 79892 125560 79898
rect 125508 79834 125560 79840
rect 125520 77897 125548 79834
rect 125658 79744 125686 80036
rect 125750 79966 125778 80036
rect 125738 79960 125790 79966
rect 125738 79902 125790 79908
rect 125842 79898 125870 80036
rect 125830 79892 125882 79898
rect 125830 79834 125882 79840
rect 125612 79716 125686 79744
rect 125934 79744 125962 80036
rect 126026 79966 126054 80036
rect 126014 79960 126066 79966
rect 126118 79937 126146 80036
rect 126210 79966 126238 80036
rect 126302 79966 126330 80036
rect 126394 79966 126422 80036
rect 126486 79966 126514 80036
rect 126198 79960 126250 79966
rect 126014 79902 126066 79908
rect 126104 79928 126160 79937
rect 126198 79902 126250 79908
rect 126290 79960 126342 79966
rect 126290 79902 126342 79908
rect 126382 79960 126434 79966
rect 126382 79902 126434 79908
rect 126474 79960 126526 79966
rect 126578 79937 126606 80036
rect 126670 79966 126698 80036
rect 126762 79971 126790 80036
rect 126658 79960 126710 79966
rect 126474 79902 126526 79908
rect 126564 79928 126620 79937
rect 126104 79863 126160 79872
rect 126658 79902 126710 79908
rect 126748 79962 126804 79971
rect 126854 79966 126882 80036
rect 126748 79897 126804 79906
rect 126842 79960 126894 79966
rect 126842 79902 126894 79908
rect 126564 79863 126620 79872
rect 126290 79824 126342 79830
rect 126164 79784 126290 79812
rect 125934 79716 126100 79744
rect 125506 77888 125562 77897
rect 125506 77823 125562 77832
rect 125612 75177 125640 79716
rect 125876 79620 125928 79626
rect 125876 79562 125928 79568
rect 125692 79484 125744 79490
rect 125692 79426 125744 79432
rect 125598 75168 125654 75177
rect 125598 75103 125654 75112
rect 125416 72412 125468 72418
rect 125416 72354 125468 72360
rect 125324 61396 125376 61402
rect 125324 61338 125376 61344
rect 125232 57248 125284 57254
rect 125232 57190 125284 57196
rect 125140 51740 125192 51746
rect 125140 51682 125192 51688
rect 124956 6248 125008 6254
rect 124956 6190 125008 6196
rect 124864 3528 124916 3534
rect 124864 3470 124916 3476
rect 125704 3466 125732 79426
rect 125782 77752 125838 77761
rect 125782 77687 125838 77696
rect 125796 4894 125824 77687
rect 125784 4888 125836 4894
rect 125784 4830 125836 4836
rect 125888 4826 125916 79562
rect 125968 78872 126020 78878
rect 125968 78814 126020 78820
rect 125980 78062 126008 78814
rect 126072 78198 126100 79716
rect 126060 78192 126112 78198
rect 126060 78134 126112 78140
rect 125968 78056 126020 78062
rect 125968 77998 126020 78004
rect 126164 77976 126192 79784
rect 126290 79766 126342 79772
rect 126704 79824 126756 79830
rect 126704 79766 126756 79772
rect 126336 79688 126388 79694
rect 126072 77948 126192 77976
rect 126256 79648 126336 79676
rect 125968 75200 126020 75206
rect 125968 75142 126020 75148
rect 125980 6186 126008 75142
rect 126072 8974 126100 77948
rect 126256 75914 126284 79648
rect 126336 79630 126388 79636
rect 126336 78192 126388 78198
rect 126336 78134 126388 78140
rect 126428 78192 126480 78198
rect 126428 78134 126480 78140
rect 126164 75886 126284 75914
rect 126164 21418 126192 75886
rect 126348 74050 126376 78134
rect 126336 74044 126388 74050
rect 126336 73986 126388 73992
rect 126440 73930 126468 78134
rect 126716 77654 126744 79766
rect 126796 79756 126848 79762
rect 126796 79698 126848 79704
rect 126704 77648 126756 77654
rect 126704 77590 126756 77596
rect 126348 73902 126468 73930
rect 126244 73228 126296 73234
rect 126244 73170 126296 73176
rect 126152 21412 126204 21418
rect 126152 21354 126204 21360
rect 126060 8968 126112 8974
rect 126060 8910 126112 8916
rect 125968 6180 126020 6186
rect 125968 6122 126020 6128
rect 125876 4820 125928 4826
rect 125876 4762 125928 4768
rect 126256 3670 126284 73170
rect 126348 18698 126376 73902
rect 126808 70394 126836 79698
rect 126946 79642 126974 80036
rect 127038 79830 127066 80036
rect 127130 79971 127158 80036
rect 127116 79962 127172 79971
rect 127116 79897 127172 79906
rect 127222 79898 127250 80036
rect 127314 79971 127342 80036
rect 127300 79962 127356 79971
rect 127210 79892 127262 79898
rect 127300 79897 127356 79906
rect 127210 79834 127262 79840
rect 127406 79830 127434 80036
rect 127498 79966 127526 80036
rect 127486 79960 127538 79966
rect 127590 79937 127618 80036
rect 127486 79902 127538 79908
rect 127576 79928 127632 79937
rect 127576 79863 127632 79872
rect 127026 79824 127078 79830
rect 127026 79766 127078 79772
rect 127394 79824 127446 79830
rect 127394 79766 127446 79772
rect 127164 79756 127216 79762
rect 127164 79698 127216 79704
rect 127256 79756 127308 79762
rect 127256 79698 127308 79704
rect 127532 79756 127584 79762
rect 127682 79744 127710 80036
rect 127774 79971 127802 80036
rect 127760 79962 127816 79971
rect 127866 79966 127894 80036
rect 127958 79966 127986 80036
rect 127760 79897 127816 79906
rect 127854 79960 127906 79966
rect 127854 79902 127906 79908
rect 127946 79960 127998 79966
rect 127946 79902 127998 79908
rect 127808 79756 127860 79762
rect 127682 79716 127756 79744
rect 127532 79698 127584 79704
rect 126900 79614 126974 79642
rect 127072 79688 127124 79694
rect 127072 79630 127124 79636
rect 126900 75206 126928 79614
rect 127084 77994 127112 79630
rect 127072 77988 127124 77994
rect 127072 77930 127124 77936
rect 127072 77308 127124 77314
rect 127072 77250 127124 77256
rect 127084 75256 127112 77250
rect 127176 76537 127204 79698
rect 127162 76528 127218 76537
rect 127162 76463 127218 76472
rect 127268 75914 127296 79698
rect 127348 79688 127400 79694
rect 127348 79630 127400 79636
rect 127360 78169 127388 79630
rect 127440 78940 127492 78946
rect 127440 78882 127492 78888
rect 127346 78160 127402 78169
rect 127346 78095 127402 78104
rect 127452 77994 127480 78882
rect 127544 78878 127572 79698
rect 127624 79484 127676 79490
rect 127624 79426 127676 79432
rect 127532 78872 127584 78878
rect 127532 78814 127584 78820
rect 127636 78112 127664 79426
rect 127728 78946 127756 79716
rect 128050 79744 128078 80036
rect 128142 79898 128170 80036
rect 128234 79966 128262 80036
rect 128222 79960 128274 79966
rect 128326 79937 128354 80036
rect 128418 79966 128446 80036
rect 128510 79966 128538 80036
rect 128406 79960 128458 79966
rect 128222 79902 128274 79908
rect 128312 79928 128368 79937
rect 128130 79892 128182 79898
rect 128406 79902 128458 79908
rect 128498 79960 128550 79966
rect 128498 79902 128550 79908
rect 128602 79898 128630 80036
rect 128694 79937 128722 80036
rect 128680 79928 128736 79937
rect 128312 79863 128368 79872
rect 128590 79892 128642 79898
rect 128130 79834 128182 79840
rect 128680 79863 128736 79872
rect 128590 79834 128642 79840
rect 128786 79830 128814 80036
rect 128878 79898 128906 80036
rect 128866 79892 128918 79898
rect 128866 79834 128918 79840
rect 128970 79830 128998 80036
rect 129062 79966 129090 80036
rect 129154 79966 129182 80036
rect 129050 79960 129102 79966
rect 129050 79902 129102 79908
rect 129142 79960 129194 79966
rect 129246 79937 129274 80036
rect 129142 79902 129194 79908
rect 129232 79928 129288 79937
rect 129338 79898 129366 80036
rect 129232 79863 129288 79872
rect 129326 79892 129378 79898
rect 129326 79834 129378 79840
rect 128774 79824 128826 79830
rect 128774 79766 128826 79772
rect 128958 79824 129010 79830
rect 128958 79766 129010 79772
rect 129188 79824 129240 79830
rect 129188 79766 129240 79772
rect 128176 79756 128228 79762
rect 128050 79716 128124 79744
rect 127808 79698 127860 79704
rect 127716 78940 127768 78946
rect 127716 78882 127768 78888
rect 127716 78804 127768 78810
rect 127716 78746 127768 78752
rect 127544 78084 127664 78112
rect 127440 77988 127492 77994
rect 127440 77930 127492 77936
rect 127438 77888 127494 77897
rect 127438 77823 127494 77832
rect 127268 75886 127388 75914
rect 127164 75472 127216 75478
rect 127164 75414 127216 75420
rect 127176 75342 127204 75414
rect 127164 75336 127216 75342
rect 127164 75278 127216 75284
rect 127256 75336 127308 75342
rect 127256 75278 127308 75284
rect 126992 75228 127112 75256
rect 126888 75200 126940 75206
rect 126888 75142 126940 75148
rect 126440 70366 126836 70394
rect 126336 18692 126388 18698
rect 126336 18634 126388 18640
rect 126244 3664 126296 3670
rect 126244 3606 126296 3612
rect 126440 3602 126468 70366
rect 126428 3596 126480 3602
rect 126428 3538 126480 3544
rect 126992 3534 127020 75228
rect 127164 75200 127216 75206
rect 127164 75142 127216 75148
rect 127072 75132 127124 75138
rect 127072 75074 127124 75080
rect 127084 4962 127112 75074
rect 127176 5098 127204 75142
rect 127268 6322 127296 75278
rect 127360 7682 127388 75886
rect 127452 75138 127480 77823
rect 127440 75132 127492 75138
rect 127440 75074 127492 75080
rect 127440 74996 127492 75002
rect 127440 74938 127492 74944
rect 127452 10334 127480 74938
rect 127544 44946 127572 78084
rect 127624 77988 127676 77994
rect 127624 77930 127676 77936
rect 127532 44940 127584 44946
rect 127532 44882 127584 44888
rect 127636 44878 127664 77930
rect 127728 75478 127756 78746
rect 127716 75472 127768 75478
rect 127716 75414 127768 75420
rect 127820 75206 127848 79698
rect 127990 79656 128046 79665
rect 127990 79591 128046 79600
rect 127900 79348 127952 79354
rect 127900 79290 127952 79296
rect 127912 79082 127940 79290
rect 127900 79076 127952 79082
rect 127900 79018 127952 79024
rect 127900 78124 127952 78130
rect 127900 78066 127952 78072
rect 127912 77314 127940 78066
rect 127900 77308 127952 77314
rect 127900 77250 127952 77256
rect 127808 75200 127860 75206
rect 127808 75142 127860 75148
rect 128004 75070 128032 79591
rect 128096 77382 128124 79716
rect 128176 79698 128228 79704
rect 128360 79756 128412 79762
rect 128360 79698 128412 79704
rect 128084 77376 128136 77382
rect 128084 77318 128136 77324
rect 128188 75914 128216 79698
rect 128266 79656 128322 79665
rect 128266 79591 128322 79600
rect 128096 75886 128216 75914
rect 128096 75342 128124 75886
rect 128084 75336 128136 75342
rect 128084 75278 128136 75284
rect 127992 75064 128044 75070
rect 127992 75006 128044 75012
rect 128280 75002 128308 79591
rect 128372 78849 128400 79698
rect 128452 79688 128504 79694
rect 128452 79630 128504 79636
rect 128544 79688 128596 79694
rect 128728 79688 128780 79694
rect 128544 79630 128596 79636
rect 128726 79656 128728 79665
rect 129096 79688 129148 79694
rect 128780 79656 128782 79665
rect 128358 78840 128414 78849
rect 128358 78775 128414 78784
rect 128360 78668 128412 78674
rect 128360 78610 128412 78616
rect 128268 74996 128320 75002
rect 128268 74938 128320 74944
rect 127624 44872 127676 44878
rect 127624 44814 127676 44820
rect 128372 10470 128400 78610
rect 128464 76673 128492 79630
rect 128556 78606 128584 79630
rect 129096 79630 129148 79636
rect 128726 79591 128782 79600
rect 128820 79620 128872 79626
rect 128820 79562 128872 79568
rect 128728 79348 128780 79354
rect 128728 79290 128780 79296
rect 128740 79150 128768 79290
rect 128728 79144 128780 79150
rect 128728 79086 128780 79092
rect 128544 78600 128596 78606
rect 128544 78542 128596 78548
rect 128544 78464 128596 78470
rect 128544 78406 128596 78412
rect 128556 76702 128584 78406
rect 128544 76696 128596 76702
rect 128450 76664 128506 76673
rect 128544 76638 128596 76644
rect 128450 76599 128506 76608
rect 128544 75336 128596 75342
rect 128544 75278 128596 75284
rect 128360 10464 128412 10470
rect 128360 10406 128412 10412
rect 127440 10328 127492 10334
rect 127440 10270 127492 10276
rect 128556 9110 128584 75278
rect 128728 75268 128780 75274
rect 128728 75210 128780 75216
rect 128636 75200 128688 75206
rect 128636 75142 128688 75148
rect 128648 9178 128676 75142
rect 128636 9172 128688 9178
rect 128636 9114 128688 9120
rect 128544 9104 128596 9110
rect 128544 9046 128596 9052
rect 128740 9042 128768 75210
rect 128832 18630 128860 79562
rect 128912 79552 128964 79558
rect 128912 79494 128964 79500
rect 128820 18624 128872 18630
rect 128820 18566 128872 18572
rect 128728 9036 128780 9042
rect 128728 8978 128780 8984
rect 127348 7676 127400 7682
rect 127348 7618 127400 7624
rect 128924 6390 128952 79494
rect 129004 79484 129056 79490
rect 129004 79426 129056 79432
rect 129016 75410 129044 79426
rect 129004 75404 129056 75410
rect 129004 75346 129056 75352
rect 129108 75274 129136 79630
rect 129200 78402 129228 79766
rect 129430 79744 129458 80036
rect 129522 79966 129550 80036
rect 129614 79966 129642 80036
rect 129510 79960 129562 79966
rect 129510 79902 129562 79908
rect 129602 79960 129654 79966
rect 129602 79902 129654 79908
rect 129706 79778 129734 80036
rect 129798 79898 129826 80036
rect 129890 79937 129918 80036
rect 129876 79928 129932 79937
rect 129786 79892 129838 79898
rect 129876 79863 129932 79872
rect 129786 79834 129838 79840
rect 129982 79830 130010 80036
rect 130074 79937 130102 80036
rect 130166 79966 130194 80036
rect 130258 79966 130286 80036
rect 130154 79960 130206 79966
rect 130060 79928 130116 79937
rect 130154 79902 130206 79908
rect 130246 79960 130298 79966
rect 130246 79902 130298 79908
rect 130060 79863 130116 79872
rect 129384 79716 129458 79744
rect 129660 79750 129734 79778
rect 129970 79824 130022 79830
rect 129970 79766 130022 79772
rect 130108 79824 130160 79830
rect 130108 79766 130160 79772
rect 129280 79688 129332 79694
rect 129280 79630 129332 79636
rect 129188 78396 129240 78402
rect 129188 78338 129240 78344
rect 129188 77784 129240 77790
rect 129188 77726 129240 77732
rect 129096 75268 129148 75274
rect 129096 75210 129148 75216
rect 129200 75154 129228 77726
rect 129108 75126 129228 75154
rect 129108 64874 129136 75126
rect 129292 70394 129320 79630
rect 129384 78810 129412 79716
rect 129556 79620 129608 79626
rect 129556 79562 129608 79568
rect 129372 78804 129424 78810
rect 129372 78746 129424 78752
rect 129370 78704 129426 78713
rect 129370 78639 129426 78648
rect 129384 75138 129412 78639
rect 129568 75206 129596 79562
rect 129660 75342 129688 79750
rect 129740 79688 129792 79694
rect 129740 79630 129792 79636
rect 130016 79688 130068 79694
rect 130016 79630 130068 79636
rect 129752 78849 129780 79630
rect 129832 79552 129884 79558
rect 129832 79494 129884 79500
rect 129738 78840 129794 78849
rect 129738 78775 129794 78784
rect 129738 77888 129794 77897
rect 129738 77823 129794 77832
rect 129752 77586 129780 77823
rect 129844 77790 129872 79494
rect 129924 79484 129976 79490
rect 129924 79426 129976 79432
rect 129832 77784 129884 77790
rect 129832 77726 129884 77732
rect 129740 77580 129792 77586
rect 129740 77522 129792 77528
rect 129648 75336 129700 75342
rect 129648 75278 129700 75284
rect 129556 75200 129608 75206
rect 129556 75142 129608 75148
rect 129740 75200 129792 75206
rect 129740 75142 129792 75148
rect 129372 75132 129424 75138
rect 129372 75074 129424 75080
rect 129016 64846 129136 64874
rect 129200 70366 129320 70394
rect 129016 9314 129044 64846
rect 129004 9308 129056 9314
rect 129004 9250 129056 9256
rect 129200 7750 129228 70366
rect 129752 16574 129780 75142
rect 129752 16546 129872 16574
rect 129188 7744 129240 7750
rect 129188 7686 129240 7692
rect 128912 6384 128964 6390
rect 128912 6326 128964 6332
rect 127256 6316 127308 6322
rect 127256 6258 127308 6264
rect 127164 5092 127216 5098
rect 127164 5034 127216 5040
rect 127072 4956 127124 4962
rect 127072 4898 127124 4904
rect 127072 3664 127124 3670
rect 127072 3606 127124 3612
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 125692 3460 125744 3466
rect 125692 3402 125744 3408
rect 127084 3346 127112 3606
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 126992 3318 127112 3346
rect 125876 3052 125928 3058
rect 125876 2994 125928 3000
rect 125888 480 125916 2994
rect 126992 480 127020 3318
rect 128188 480 128216 3470
rect 129384 480 129412 3538
rect 129844 3482 129872 16546
rect 129936 5166 129964 79426
rect 130028 78713 130056 79630
rect 130014 78704 130070 78713
rect 130014 78639 130070 78648
rect 130016 75268 130068 75274
rect 130016 75210 130068 75216
rect 130028 6458 130056 75210
rect 130120 9246 130148 79766
rect 130350 79744 130378 80036
rect 130442 79898 130470 80036
rect 130430 79892 130482 79898
rect 130430 79834 130482 79840
rect 130534 79744 130562 80036
rect 130626 79898 130654 80036
rect 130718 79966 130746 80036
rect 130706 79960 130758 79966
rect 130706 79902 130758 79908
rect 130810 79898 130838 80036
rect 130902 79966 130930 80036
rect 130994 79966 131022 80036
rect 131086 79966 131114 80036
rect 131178 79971 131206 80036
rect 130890 79960 130942 79966
rect 130890 79902 130942 79908
rect 130982 79960 131034 79966
rect 130982 79902 131034 79908
rect 131074 79960 131126 79966
rect 131074 79902 131126 79908
rect 131164 79962 131220 79971
rect 131270 79966 131298 80036
rect 130614 79892 130666 79898
rect 130614 79834 130666 79840
rect 130798 79892 130850 79898
rect 131164 79897 131220 79906
rect 131258 79960 131310 79966
rect 131362 79937 131390 80036
rect 131454 79966 131482 80036
rect 131546 79966 131574 80036
rect 131638 79966 131666 80036
rect 131442 79960 131494 79966
rect 131258 79902 131310 79908
rect 131348 79928 131404 79937
rect 131442 79902 131494 79908
rect 131534 79960 131586 79966
rect 131534 79902 131586 79908
rect 131626 79960 131678 79966
rect 131626 79902 131678 79908
rect 131348 79863 131404 79872
rect 130798 79834 130850 79840
rect 130890 79824 130942 79830
rect 130350 79716 130424 79744
rect 130292 79416 130344 79422
rect 130292 79358 130344 79364
rect 130200 77988 130252 77994
rect 130200 77930 130252 77936
rect 130212 73914 130240 77930
rect 130200 73908 130252 73914
rect 130200 73850 130252 73856
rect 130304 70394 130332 79358
rect 130396 77994 130424 79716
rect 130488 79716 130562 79744
rect 130810 79772 130890 79778
rect 130810 79766 130942 79772
rect 131580 79824 131632 79830
rect 131730 79812 131758 80036
rect 131822 79966 131850 80036
rect 131810 79960 131862 79966
rect 131810 79902 131862 79908
rect 131730 79784 131804 79812
rect 131580 79766 131632 79772
rect 130810 79750 130930 79766
rect 131304 79756 131356 79762
rect 130488 78198 130516 79716
rect 130660 79688 130712 79694
rect 130810 79676 130838 79750
rect 131304 79698 131356 79704
rect 130936 79688 130988 79694
rect 130810 79648 130884 79676
rect 130660 79630 130712 79636
rect 130568 79620 130620 79626
rect 130568 79562 130620 79568
rect 130476 78192 130528 78198
rect 130476 78134 130528 78140
rect 130384 77988 130436 77994
rect 130384 77930 130436 77936
rect 130476 77308 130528 77314
rect 130476 77250 130528 77256
rect 130488 75206 130516 77250
rect 130476 75200 130528 75206
rect 130476 75142 130528 75148
rect 130476 74520 130528 74526
rect 130382 74488 130438 74497
rect 130476 74462 130528 74468
rect 130382 74423 130438 74432
rect 130212 70366 130332 70394
rect 130212 45014 130240 70366
rect 130200 45008 130252 45014
rect 130200 44950 130252 44956
rect 130108 9240 130160 9246
rect 130108 9182 130160 9188
rect 130396 6914 130424 74423
rect 130304 6886 130424 6914
rect 130016 6452 130068 6458
rect 130016 6394 130068 6400
rect 129924 5160 129976 5166
rect 129924 5102 129976 5108
rect 130304 3670 130332 6886
rect 130292 3664 130344 3670
rect 130292 3606 130344 3612
rect 130488 3602 130516 74462
rect 130580 16574 130608 79562
rect 130672 75274 130700 79630
rect 130660 75268 130712 75274
rect 130660 75210 130712 75216
rect 130856 73234 130884 79648
rect 130936 79630 130988 79636
rect 131212 79688 131264 79694
rect 131212 79630 131264 79636
rect 130948 76634 130976 79630
rect 131120 79620 131172 79626
rect 131120 79562 131172 79568
rect 131132 77294 131160 79562
rect 131224 78713 131252 79630
rect 131210 78704 131266 78713
rect 131210 78639 131266 78648
rect 131316 77994 131344 79698
rect 131488 79620 131540 79626
rect 131488 79562 131540 79568
rect 131304 77988 131356 77994
rect 131304 77930 131356 77936
rect 131304 77784 131356 77790
rect 131304 77726 131356 77732
rect 131132 77266 131252 77294
rect 131224 76770 131252 77266
rect 131212 76764 131264 76770
rect 131212 76706 131264 76712
rect 130936 76628 130988 76634
rect 130936 76570 130988 76576
rect 131212 75200 131264 75206
rect 131212 75142 131264 75148
rect 130844 73228 130896 73234
rect 130844 73170 130896 73176
rect 130580 16546 130700 16574
rect 130672 3738 130700 16546
rect 131224 4078 131252 75142
rect 131212 4072 131264 4078
rect 131212 4014 131264 4020
rect 131316 3874 131344 77726
rect 131396 75268 131448 75274
rect 131396 75210 131448 75216
rect 131408 6594 131436 75210
rect 131396 6588 131448 6594
rect 131396 6530 131448 6536
rect 131500 6526 131528 79562
rect 131592 78674 131620 79766
rect 131580 78668 131632 78674
rect 131580 78610 131632 78616
rect 131580 78260 131632 78266
rect 131580 78202 131632 78208
rect 131592 7818 131620 78202
rect 131670 78160 131726 78169
rect 131670 78095 131726 78104
rect 131684 10606 131712 78095
rect 131776 77790 131804 79784
rect 131914 79744 131942 80036
rect 132006 79830 132034 80036
rect 132098 79898 132126 80036
rect 132190 79971 132218 80036
rect 132176 79962 132232 79971
rect 132282 79966 132310 80036
rect 132374 79966 132402 80036
rect 132466 79966 132494 80036
rect 132558 79971 132586 80036
rect 132086 79892 132138 79898
rect 132176 79897 132232 79906
rect 132270 79960 132322 79966
rect 132270 79902 132322 79908
rect 132362 79960 132414 79966
rect 132362 79902 132414 79908
rect 132454 79960 132506 79966
rect 132454 79902 132506 79908
rect 132544 79962 132600 79971
rect 132544 79897 132600 79906
rect 132650 79898 132678 80036
rect 132742 79898 132770 80036
rect 132834 79966 132862 80036
rect 132822 79960 132874 79966
rect 132822 79902 132874 79908
rect 132086 79834 132138 79840
rect 132638 79892 132690 79898
rect 132638 79834 132690 79840
rect 132730 79892 132782 79898
rect 132730 79834 132782 79840
rect 131994 79824 132046 79830
rect 131994 79766 132046 79772
rect 132774 79792 132830 79801
rect 131868 79716 131942 79744
rect 132224 79756 132276 79762
rect 131764 77784 131816 77790
rect 131764 77726 131816 77732
rect 131868 70394 131896 79716
rect 132224 79698 132276 79704
rect 132592 79756 132644 79762
rect 132926 79744 132954 80036
rect 133018 79971 133046 80036
rect 133004 79962 133060 79971
rect 133004 79897 133060 79906
rect 133110 79898 133138 80036
rect 133202 79966 133230 80036
rect 133190 79960 133242 79966
rect 133190 79902 133242 79908
rect 133098 79892 133150 79898
rect 133098 79834 133150 79840
rect 133294 79778 133322 80036
rect 132774 79727 132830 79736
rect 132592 79698 132644 79704
rect 132040 79688 132092 79694
rect 132040 79630 132092 79636
rect 132132 79688 132184 79694
rect 132132 79630 132184 79636
rect 131948 79620 132000 79626
rect 131948 79562 132000 79568
rect 131960 75274 131988 79562
rect 132052 78112 132080 79630
rect 132144 78266 132172 79630
rect 132132 78260 132184 78266
rect 132132 78202 132184 78208
rect 132052 78084 132172 78112
rect 132040 77988 132092 77994
rect 132040 77930 132092 77936
rect 132052 75614 132080 77930
rect 132040 75608 132092 75614
rect 132040 75550 132092 75556
rect 131948 75268 132000 75274
rect 131948 75210 132000 75216
rect 132144 75206 132172 78084
rect 132132 75200 132184 75206
rect 132132 75142 132184 75148
rect 132236 70394 132264 79698
rect 132316 79688 132368 79694
rect 132316 79630 132368 79636
rect 132328 77042 132356 79630
rect 132604 78033 132632 79698
rect 132684 79688 132736 79694
rect 132682 79656 132684 79665
rect 132736 79656 132738 79665
rect 132682 79591 132738 79600
rect 132684 79552 132736 79558
rect 132684 79494 132736 79500
rect 132590 78024 132646 78033
rect 132590 77959 132646 77968
rect 132316 77036 132368 77042
rect 132316 76978 132368 76984
rect 132696 76838 132724 79494
rect 132788 78062 132816 79727
rect 132880 79716 132954 79744
rect 133144 79756 133196 79762
rect 132880 78470 132908 79716
rect 133144 79698 133196 79704
rect 133248 79750 133322 79778
rect 133386 79778 133414 80036
rect 133478 79898 133506 80036
rect 133466 79892 133518 79898
rect 133466 79834 133518 79840
rect 133570 79778 133598 80036
rect 133662 79966 133690 80036
rect 133650 79960 133702 79966
rect 133650 79902 133702 79908
rect 133386 79750 133460 79778
rect 133052 79620 133104 79626
rect 133052 79562 133104 79568
rect 132868 78464 132920 78470
rect 132868 78406 132920 78412
rect 132776 78056 132828 78062
rect 133064 78010 133092 79562
rect 132776 77998 132828 78004
rect 132880 77982 133092 78010
rect 132684 76832 132736 76838
rect 132684 76774 132736 76780
rect 132684 75336 132736 75342
rect 132684 75278 132736 75284
rect 131776 70366 131896 70394
rect 132144 70366 132264 70394
rect 131672 10600 131724 10606
rect 131672 10542 131724 10548
rect 131776 10538 131804 70366
rect 132144 64874 132172 70366
rect 131868 64846 132172 64874
rect 131764 10532 131816 10538
rect 131764 10474 131816 10480
rect 131580 7812 131632 7818
rect 131580 7754 131632 7760
rect 131488 6520 131540 6526
rect 131488 6462 131540 6468
rect 131868 4010 131896 64846
rect 132696 6662 132724 75278
rect 132776 75200 132828 75206
rect 132776 75142 132828 75148
rect 132788 7954 132816 75142
rect 132776 7948 132828 7954
rect 132776 7890 132828 7896
rect 132880 7886 132908 77982
rect 132960 76492 133012 76498
rect 132960 76434 133012 76440
rect 132972 10402 133000 76434
rect 133052 75268 133104 75274
rect 133052 75210 133104 75216
rect 133064 11762 133092 75210
rect 133156 72486 133184 79698
rect 133248 76498 133276 79750
rect 133432 79676 133460 79750
rect 133386 79648 133460 79676
rect 133524 79750 133598 79778
rect 133386 79642 133414 79648
rect 133340 79614 133414 79642
rect 133236 76492 133288 76498
rect 133236 76434 133288 76440
rect 133144 72480 133196 72486
rect 133144 72422 133196 72428
rect 133340 70394 133368 79614
rect 133524 79608 133552 79750
rect 133754 79744 133782 80036
rect 133708 79716 133782 79744
rect 133604 79688 133656 79694
rect 133604 79630 133656 79636
rect 133478 79580 133552 79608
rect 133478 79540 133506 79580
rect 133432 79512 133506 79540
rect 133432 77926 133460 79512
rect 133512 79416 133564 79422
rect 133512 79358 133564 79364
rect 133420 77920 133472 77926
rect 133420 77862 133472 77868
rect 133156 70366 133368 70394
rect 133052 11756 133104 11762
rect 133052 11698 133104 11704
rect 132960 10396 133012 10402
rect 132960 10338 133012 10344
rect 132868 7880 132920 7886
rect 132868 7822 132920 7828
rect 132684 6656 132736 6662
rect 132684 6598 132736 6604
rect 133156 5302 133184 70366
rect 133524 64874 133552 79358
rect 133616 75342 133644 79630
rect 133604 75336 133656 75342
rect 133604 75278 133656 75284
rect 133708 75206 133736 79716
rect 133846 79676 133874 80036
rect 133938 79937 133966 80036
rect 134030 79966 134058 80036
rect 134018 79960 134070 79966
rect 133924 79928 133980 79937
rect 134018 79902 134070 79908
rect 133924 79863 133980 79872
rect 134122 79830 134150 80036
rect 134214 79898 134242 80036
rect 134306 79937 134334 80036
rect 134292 79928 134348 79937
rect 134202 79892 134254 79898
rect 134398 79898 134426 80036
rect 134490 79971 134518 80036
rect 134476 79962 134532 79971
rect 134582 79966 134610 80036
rect 134292 79863 134348 79872
rect 134386 79892 134438 79898
rect 134476 79897 134532 79906
rect 134570 79960 134622 79966
rect 134570 79902 134622 79908
rect 134202 79834 134254 79840
rect 134386 79834 134438 79840
rect 133972 79824 134024 79830
rect 133972 79766 134024 79772
rect 134110 79824 134162 79830
rect 134110 79766 134162 79772
rect 134430 79792 134486 79801
rect 133800 79648 133874 79676
rect 133800 75274 133828 79648
rect 133880 78192 133932 78198
rect 133880 78134 133932 78140
rect 133788 75268 133840 75274
rect 133788 75210 133840 75216
rect 133696 75200 133748 75206
rect 133696 75142 133748 75148
rect 133340 64846 133552 64874
rect 133144 5296 133196 5302
rect 133144 5238 133196 5244
rect 133340 5234 133368 64846
rect 133328 5228 133380 5234
rect 133328 5170 133380 5176
rect 131856 4004 131908 4010
rect 131856 3946 131908 3952
rect 131304 3868 131356 3874
rect 131304 3810 131356 3816
rect 130660 3732 130712 3738
rect 130660 3674 130712 3680
rect 130476 3596 130528 3602
rect 130476 3538 130528 3544
rect 129844 3454 130608 3482
rect 130580 480 130608 3454
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 131776 480 131804 3402
rect 132960 3120 133012 3126
rect 132960 3062 133012 3068
rect 132972 480 133000 3062
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 78134
rect 133984 78033 134012 79766
rect 134674 79778 134702 80036
rect 134766 79937 134794 80036
rect 134858 79966 134886 80036
rect 134950 79971 134978 80036
rect 134846 79960 134898 79966
rect 134752 79928 134808 79937
rect 134846 79902 134898 79908
rect 134936 79962 134992 79971
rect 134936 79897 134992 79906
rect 135042 79898 135070 80036
rect 134752 79863 134808 79872
rect 135030 79892 135082 79898
rect 135030 79834 135082 79840
rect 134982 79792 135038 79801
rect 134430 79727 134486 79736
rect 134524 79756 134576 79762
rect 134338 79656 134394 79665
rect 134064 79620 134116 79626
rect 134064 79562 134116 79568
rect 134248 79620 134300 79626
rect 134338 79591 134394 79600
rect 134248 79562 134300 79568
rect 134076 78713 134104 79562
rect 134156 79552 134208 79558
rect 134156 79494 134208 79500
rect 134062 78704 134118 78713
rect 134062 78639 134118 78648
rect 134064 78260 134116 78266
rect 134064 78202 134116 78208
rect 133970 78024 134026 78033
rect 133970 77959 134026 77968
rect 134076 77518 134104 78202
rect 134064 77512 134116 77518
rect 134064 77454 134116 77460
rect 134168 75914 134196 79494
rect 134260 78266 134288 79562
rect 134248 78260 134300 78266
rect 134248 78202 134300 78208
rect 134248 78056 134300 78062
rect 134248 77998 134300 78004
rect 134076 75886 134196 75914
rect 134076 5370 134104 75886
rect 134156 75268 134208 75274
rect 134156 75210 134208 75216
rect 134168 8022 134196 75210
rect 134260 11830 134288 77998
rect 134352 76809 134380 79591
rect 134444 78334 134472 79727
rect 134674 79750 134932 79778
rect 134524 79698 134576 79704
rect 134432 78328 134484 78334
rect 134432 78270 134484 78276
rect 134432 77988 134484 77994
rect 134432 77930 134484 77936
rect 134338 76800 134394 76809
rect 134338 76735 134394 76744
rect 134444 73982 134472 77930
rect 134536 75274 134564 79698
rect 134616 79688 134668 79694
rect 134616 79630 134668 79636
rect 134708 79688 134760 79694
rect 134708 79630 134760 79636
rect 134798 79656 134854 79665
rect 134628 76906 134656 79630
rect 134616 76900 134668 76906
rect 134616 76842 134668 76848
rect 134720 75914 134748 79630
rect 134798 79591 134854 79600
rect 134812 77994 134840 79591
rect 134904 78062 134932 79750
rect 134982 79727 135038 79736
rect 135134 79744 135162 80036
rect 135226 79966 135254 80036
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 135318 79898 135346 80036
rect 135410 79937 135438 80036
rect 135502 79966 135530 80036
rect 135594 79966 135622 80036
rect 135490 79960 135542 79966
rect 135396 79928 135452 79937
rect 135306 79892 135358 79898
rect 135490 79902 135542 79908
rect 135582 79960 135634 79966
rect 135686 79937 135714 80036
rect 135582 79902 135634 79908
rect 135672 79928 135728 79937
rect 135396 79863 135452 79872
rect 135672 79863 135728 79872
rect 135306 79834 135358 79840
rect 135778 79830 135806 80036
rect 135870 79966 135898 80036
rect 135858 79960 135910 79966
rect 135858 79902 135910 79908
rect 135766 79824 135818 79830
rect 135766 79766 135818 79772
rect 135962 79778 135990 80036
rect 136054 79898 136082 80036
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 136146 79778 136174 80036
rect 136238 79966 136266 80036
rect 136330 79966 136358 80036
rect 136422 79966 136450 80036
rect 136514 79971 136542 80036
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 136410 79960 136462 79966
rect 136410 79902 136462 79908
rect 136500 79962 136556 79971
rect 136606 79966 136634 80036
rect 136500 79897 136556 79906
rect 136594 79960 136646 79966
rect 136594 79902 136646 79908
rect 136698 79830 136726 80036
rect 136790 79971 136818 80036
rect 136776 79962 136832 79971
rect 136776 79897 136832 79906
rect 136686 79824 136738 79830
rect 135352 79756 135404 79762
rect 134892 78056 134944 78062
rect 134892 77998 134944 78004
rect 134800 77988 134852 77994
rect 134800 77930 134852 77936
rect 134996 77450 135024 79727
rect 135134 79716 135208 79744
rect 135076 79620 135128 79626
rect 135076 79562 135128 79568
rect 134984 77444 135036 77450
rect 134984 77386 135036 77392
rect 134628 75886 134748 75914
rect 134628 75546 134656 75886
rect 134616 75540 134668 75546
rect 134616 75482 134668 75488
rect 134524 75268 134576 75274
rect 134524 75210 134576 75216
rect 134432 73976 134484 73982
rect 134432 73918 134484 73924
rect 135088 70394 135116 79562
rect 135180 76974 135208 79716
rect 135352 79698 135404 79704
rect 135444 79756 135496 79762
rect 135962 79750 136036 79778
rect 135444 79698 135496 79704
rect 135260 79620 135312 79626
rect 135260 79562 135312 79568
rect 135168 76968 135220 76974
rect 135168 76910 135220 76916
rect 135168 76764 135220 76770
rect 135168 76706 135220 76712
rect 134904 70366 135116 70394
rect 134904 64874 134932 70366
rect 134536 64846 134932 64874
rect 134248 11824 134300 11830
rect 134248 11766 134300 11772
rect 134156 8016 134208 8022
rect 134156 7958 134208 7964
rect 134064 5364 134116 5370
rect 134064 5306 134116 5312
rect 134536 3942 134564 64846
rect 134524 3936 134576 3942
rect 134524 3878 134576 3884
rect 135180 3738 135208 76706
rect 135272 74526 135300 79562
rect 135364 77858 135392 79698
rect 135456 78130 135484 79698
rect 135720 79688 135772 79694
rect 135904 79688 135956 79694
rect 135720 79630 135772 79636
rect 135810 79656 135866 79665
rect 135628 79552 135680 79558
rect 135628 79494 135680 79500
rect 135536 78668 135588 78674
rect 135536 78610 135588 78616
rect 135444 78124 135496 78130
rect 135444 78066 135496 78072
rect 135352 77852 135404 77858
rect 135352 77794 135404 77800
rect 135352 75336 135404 75342
rect 135352 75278 135404 75284
rect 135260 74520 135312 74526
rect 135260 74462 135312 74468
rect 135364 6914 135392 75278
rect 135444 75132 135496 75138
rect 135444 75074 135496 75080
rect 135272 6886 135392 6914
rect 135168 3732 135220 3738
rect 135168 3674 135220 3680
rect 135272 480 135300 6886
rect 135456 3602 135484 75074
rect 135444 3596 135496 3602
rect 135444 3538 135496 3544
rect 135548 3126 135576 78610
rect 135640 75342 135668 79494
rect 135732 75914 135760 79630
rect 135904 79630 135956 79636
rect 135810 79591 135866 79600
rect 135824 77314 135852 79591
rect 135916 78674 135944 79630
rect 135904 78668 135956 78674
rect 135904 78610 135956 78616
rect 136008 78198 136036 79750
rect 136100 79750 136174 79778
rect 136454 79792 136510 79801
rect 136364 79756 136416 79762
rect 135996 78192 136048 78198
rect 135996 78134 136048 78140
rect 135996 78056 136048 78062
rect 135996 77998 136048 78004
rect 135812 77308 135864 77314
rect 135812 77250 135864 77256
rect 135732 75886 135944 75914
rect 135628 75336 135680 75342
rect 135628 75278 135680 75284
rect 135812 75336 135864 75342
rect 135812 75278 135864 75284
rect 135720 75268 135772 75274
rect 135720 75210 135772 75216
rect 135628 75200 135680 75206
rect 135628 75142 135680 75148
rect 135536 3120 135588 3126
rect 135536 3062 135588 3068
rect 135640 3058 135668 75142
rect 135732 3534 135760 75210
rect 135720 3528 135772 3534
rect 135720 3470 135772 3476
rect 135824 3194 135852 75278
rect 135916 3466 135944 75886
rect 136008 75206 136036 77998
rect 135996 75200 136048 75206
rect 135996 75142 136048 75148
rect 136100 70394 136128 79750
rect 136686 79766 136738 79772
rect 136882 79778 136910 80036
rect 136974 79971 137002 80036
rect 136960 79962 137016 79971
rect 137066 79966 137094 80036
rect 136960 79897 137016 79906
rect 137054 79960 137106 79966
rect 137054 79902 137106 79908
rect 137006 79792 137062 79801
rect 136882 79750 136956 79778
rect 136454 79727 136510 79736
rect 136364 79698 136416 79704
rect 136180 79688 136232 79694
rect 136180 79630 136232 79636
rect 136272 79688 136324 79694
rect 136272 79630 136324 79636
rect 136192 78062 136220 79630
rect 136180 78056 136232 78062
rect 136180 77998 136232 78004
rect 136284 75274 136312 79630
rect 136272 75268 136324 75274
rect 136272 75210 136324 75216
rect 136376 75138 136404 79698
rect 136468 75342 136496 79727
rect 136824 79688 136876 79694
rect 136638 79656 136694 79665
rect 136638 79591 136694 79600
rect 136744 79648 136824 79676
rect 136652 75914 136680 79591
rect 136560 75886 136680 75914
rect 136456 75336 136508 75342
rect 136456 75278 136508 75284
rect 136364 75132 136416 75138
rect 136364 75074 136416 75080
rect 136008 70366 136128 70394
rect 136008 16574 136036 70366
rect 136008 16546 136496 16574
rect 135904 3460 135956 3466
rect 135904 3402 135956 3408
rect 135812 3188 135864 3194
rect 135812 3130 135864 3136
rect 135628 3052 135680 3058
rect 135628 2994 135680 3000
rect 136468 480 136496 16546
rect 136560 3670 136588 75886
rect 136548 3664 136600 3670
rect 136548 3606 136600 3612
rect 136744 3126 136772 79648
rect 136824 79630 136876 79636
rect 136824 79552 136876 79558
rect 136824 79494 136876 79500
rect 136836 78849 136864 79494
rect 136822 78840 136878 78849
rect 136822 78775 136878 78784
rect 136824 78668 136876 78674
rect 136824 78610 136876 78616
rect 136836 4078 136864 78610
rect 136928 5030 136956 79750
rect 137006 79727 137062 79736
rect 137158 79744 137186 80036
rect 137250 79937 137278 80036
rect 137236 79928 137292 79937
rect 137342 79898 137370 80036
rect 137434 79971 137462 80036
rect 137420 79962 137476 79971
rect 137236 79863 137292 79872
rect 137330 79892 137382 79898
rect 137420 79897 137476 79906
rect 137330 79834 137382 79840
rect 137526 79744 137554 80036
rect 137618 79966 137646 80036
rect 137710 79966 137738 80036
rect 137606 79960 137658 79966
rect 137606 79902 137658 79908
rect 137698 79960 137750 79966
rect 137698 79902 137750 79908
rect 137802 79898 137830 80036
rect 137790 79892 137842 79898
rect 137790 79834 137842 79840
rect 137894 79812 137922 80036
rect 137986 79966 138014 80036
rect 137974 79960 138026 79966
rect 138078 79937 138106 80036
rect 137974 79902 138026 79908
rect 138064 79928 138120 79937
rect 138064 79863 138120 79872
rect 138170 79812 138198 80036
rect 138262 79966 138290 80036
rect 138354 79966 138382 80036
rect 138250 79960 138302 79966
rect 138250 79902 138302 79908
rect 138342 79960 138394 79966
rect 138342 79902 138394 79908
rect 137894 79801 137968 79812
rect 137894 79792 137982 79801
rect 137894 79784 137926 79792
rect 137020 78690 137048 79727
rect 137158 79716 137232 79744
rect 137100 79076 137152 79082
rect 137100 79018 137152 79024
rect 137112 78946 137140 79018
rect 137100 78940 137152 78946
rect 137100 78882 137152 78888
rect 137020 78662 137140 78690
rect 137008 78600 137060 78606
rect 137008 78542 137060 78548
rect 137020 6322 137048 78542
rect 137112 75410 137140 78662
rect 137204 78606 137232 79716
rect 137480 79716 137554 79744
rect 138170 79784 138244 79812
rect 137926 79727 137982 79736
rect 137284 79688 137336 79694
rect 137284 79630 137336 79636
rect 137374 79656 137430 79665
rect 137192 78600 137244 78606
rect 137192 78542 137244 78548
rect 137100 75404 137152 75410
rect 137100 75346 137152 75352
rect 137100 75268 137152 75274
rect 137100 75210 137152 75216
rect 137008 6316 137060 6322
rect 137008 6258 137060 6264
rect 137112 6254 137140 75210
rect 137296 70514 137324 79630
rect 137374 79591 137430 79600
rect 137388 78674 137416 79591
rect 137376 78668 137428 78674
rect 137376 78610 137428 78616
rect 137480 75274 137508 79716
rect 137926 79656 137982 79665
rect 137926 79591 137982 79600
rect 138112 79620 138164 79626
rect 137652 79552 137704 79558
rect 137652 79494 137704 79500
rect 137744 79552 137796 79558
rect 137744 79494 137796 79500
rect 137664 77294 137692 79494
rect 137572 77266 137692 77294
rect 137468 75268 137520 75274
rect 137468 75210 137520 75216
rect 137572 73574 137600 77266
rect 137756 75914 137784 79494
rect 137940 76702 137968 79591
rect 138112 79562 138164 79568
rect 138124 78849 138152 79562
rect 138110 78840 138166 78849
rect 138110 78775 138166 78784
rect 138018 78704 138074 78713
rect 138018 78639 138074 78648
rect 138112 78668 138164 78674
rect 138032 76770 138060 78639
rect 138112 78610 138164 78616
rect 138020 76764 138072 76770
rect 138020 76706 138072 76712
rect 137928 76696 137980 76702
rect 137928 76638 137980 76644
rect 137664 75886 137784 75914
rect 137560 73568 137612 73574
rect 137560 73510 137612 73516
rect 137284 70508 137336 70514
rect 137284 70450 137336 70456
rect 137664 70394 137692 75886
rect 137744 75404 137796 75410
rect 137744 75346 137796 75352
rect 137204 70366 137692 70394
rect 137100 6248 137152 6254
rect 137100 6190 137152 6196
rect 137204 6186 137232 70366
rect 137192 6180 137244 6186
rect 137192 6122 137244 6128
rect 136916 5024 136968 5030
rect 136916 4966 136968 4972
rect 136824 4072 136876 4078
rect 136824 4014 136876 4020
rect 137756 3262 137784 75346
rect 138124 5234 138152 78610
rect 138112 5228 138164 5234
rect 138112 5170 138164 5176
rect 138216 4826 138244 79784
rect 138446 79778 138474 80036
rect 138538 79966 138566 80036
rect 138630 79966 138658 80036
rect 138722 79966 138750 80036
rect 138526 79960 138578 79966
rect 138526 79902 138578 79908
rect 138618 79960 138670 79966
rect 138618 79902 138670 79908
rect 138710 79960 138762 79966
rect 138710 79902 138762 79908
rect 138814 79898 138842 80036
rect 138906 79898 138934 80036
rect 138998 79966 139026 80036
rect 139090 79971 139118 80036
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 139076 79962 139132 79971
rect 139182 79966 139210 80036
rect 138802 79892 138854 79898
rect 138802 79834 138854 79840
rect 138894 79892 138946 79898
rect 139076 79897 139132 79906
rect 139170 79960 139222 79966
rect 139170 79902 139222 79908
rect 138894 79834 138946 79840
rect 139124 79824 139176 79830
rect 138446 79750 138612 79778
rect 139124 79766 139176 79772
rect 138388 79688 138440 79694
rect 138388 79630 138440 79636
rect 138480 79688 138532 79694
rect 138480 79630 138532 79636
rect 138296 79620 138348 79626
rect 138296 79562 138348 79568
rect 138308 75274 138336 79562
rect 138400 78334 138428 79630
rect 138388 78328 138440 78334
rect 138388 78270 138440 78276
rect 138492 75914 138520 79630
rect 138584 78674 138612 79750
rect 138664 79756 138716 79762
rect 138664 79698 138716 79704
rect 138756 79756 138808 79762
rect 138756 79698 138808 79704
rect 138940 79756 138992 79762
rect 138940 79698 138992 79704
rect 139032 79756 139084 79762
rect 139032 79698 139084 79704
rect 138572 78668 138624 78674
rect 138572 78610 138624 78616
rect 138676 78554 138704 79698
rect 138400 75886 138520 75914
rect 138584 78526 138704 78554
rect 138296 75268 138348 75274
rect 138296 75210 138348 75216
rect 138296 75132 138348 75138
rect 138296 75074 138348 75080
rect 138308 4894 138336 75074
rect 138400 4962 138428 75886
rect 138480 75268 138532 75274
rect 138480 75210 138532 75216
rect 138492 61402 138520 75210
rect 138584 75138 138612 78526
rect 138768 78418 138796 79698
rect 138848 79484 138900 79490
rect 138848 79426 138900 79432
rect 138676 78390 138796 78418
rect 138572 75132 138624 75138
rect 138572 75074 138624 75080
rect 138676 70394 138704 78390
rect 138756 78328 138808 78334
rect 138756 78270 138808 78276
rect 138768 74526 138796 78270
rect 138756 74520 138808 74526
rect 138756 74462 138808 74468
rect 138584 70366 138704 70394
rect 138756 70440 138808 70446
rect 138756 70382 138808 70388
rect 138584 67590 138612 70366
rect 138572 67584 138624 67590
rect 138572 67526 138624 67532
rect 138480 61396 138532 61402
rect 138480 61338 138532 61344
rect 138388 4956 138440 4962
rect 138388 4898 138440 4904
rect 138296 4888 138348 4894
rect 138296 4830 138348 4836
rect 138204 4820 138256 4826
rect 138204 4762 138256 4768
rect 138768 3874 138796 70382
rect 138860 4146 138888 79426
rect 138952 78606 138980 79698
rect 139044 79665 139072 79698
rect 139030 79656 139086 79665
rect 139030 79591 139086 79600
rect 139032 79552 139084 79558
rect 139032 79494 139084 79500
rect 138940 78600 138992 78606
rect 138940 78542 138992 78548
rect 138848 4140 138900 4146
rect 138848 4082 138900 4088
rect 138756 3868 138808 3874
rect 138756 3810 138808 3816
rect 138848 3528 138900 3534
rect 138848 3470 138900 3476
rect 137744 3256 137796 3262
rect 137744 3198 137796 3204
rect 136732 3120 136784 3126
rect 136732 3062 136784 3068
rect 137652 3052 137704 3058
rect 137652 2994 137704 3000
rect 137664 480 137692 2994
rect 138860 480 138888 3470
rect 139044 3330 139072 79494
rect 139136 78713 139164 79766
rect 139274 79642 139302 80036
rect 139366 79835 139394 80036
rect 139458 79971 139486 80036
rect 139444 79962 139500 79971
rect 139444 79897 139500 79906
rect 139550 79898 139578 80036
rect 139642 79966 139670 80036
rect 139734 79966 139762 80036
rect 139826 79966 139854 80036
rect 139918 79966 139946 80036
rect 140010 79966 140038 80036
rect 139630 79960 139682 79966
rect 139630 79902 139682 79908
rect 139722 79960 139774 79966
rect 139722 79902 139774 79908
rect 139814 79960 139866 79966
rect 139814 79902 139866 79908
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 139998 79960 140050 79966
rect 139998 79902 140050 79908
rect 140102 79903 140130 80036
rect 140194 79966 140222 80036
rect 140286 79966 140314 80036
rect 140378 79966 140406 80036
rect 140470 79966 140498 80036
rect 140182 79960 140234 79966
rect 139538 79892 139590 79898
rect 139352 79826 139408 79835
rect 139538 79834 139590 79840
rect 140088 79894 140144 79903
rect 140182 79902 140234 79908
rect 140274 79960 140326 79966
rect 140274 79902 140326 79908
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140458 79960 140510 79966
rect 140458 79902 140510 79908
rect 140088 79829 140144 79838
rect 140228 79824 140280 79830
rect 139352 79761 139408 79770
rect 139950 79792 140006 79801
rect 139584 79756 139636 79762
rect 139584 79698 139636 79704
rect 139676 79756 139728 79762
rect 139676 79698 139728 79704
rect 139860 79756 139912 79762
rect 140228 79766 140280 79772
rect 140412 79824 140464 79830
rect 140562 79812 140590 80036
rect 140412 79766 140464 79772
rect 140516 79784 140590 79812
rect 139950 79727 140006 79736
rect 140136 79756 140188 79762
rect 139860 79698 139912 79704
rect 139596 79665 139624 79698
rect 139582 79656 139638 79665
rect 139274 79614 139348 79642
rect 139122 78704 139178 78713
rect 139122 78639 139178 78648
rect 139124 78600 139176 78606
rect 139124 78542 139176 78548
rect 139136 71534 139164 78542
rect 139320 76362 139348 79614
rect 139582 79591 139638 79600
rect 139584 79552 139636 79558
rect 139584 79494 139636 79500
rect 139308 76356 139360 76362
rect 139308 76298 139360 76304
rect 139398 75984 139454 75993
rect 139398 75919 139454 75928
rect 139124 71528 139176 71534
rect 139124 71470 139176 71476
rect 139412 6866 139440 75919
rect 139596 75914 139624 79494
rect 139688 77994 139716 79698
rect 139768 79688 139820 79694
rect 139768 79630 139820 79636
rect 139676 77988 139728 77994
rect 139676 77930 139728 77936
rect 139504 75886 139624 75914
rect 139676 75948 139728 75954
rect 139676 75890 139728 75896
rect 139504 11558 139532 75886
rect 139584 75676 139636 75682
rect 139584 75618 139636 75624
rect 139596 14346 139624 75618
rect 139688 27198 139716 75890
rect 139780 27334 139808 79630
rect 139768 27328 139820 27334
rect 139768 27270 139820 27276
rect 139872 27266 139900 79698
rect 139964 78334 139992 79727
rect 140136 79698 140188 79704
rect 140042 79656 140098 79665
rect 140042 79591 140098 79600
rect 139952 78328 140004 78334
rect 139952 78270 140004 78276
rect 140056 75954 140084 79591
rect 140044 75948 140096 75954
rect 140044 75890 140096 75896
rect 139952 75744 140004 75750
rect 139952 75686 140004 75692
rect 139964 67114 139992 75686
rect 140148 75682 140176 79698
rect 140240 75750 140268 79766
rect 140320 79688 140372 79694
rect 140320 79630 140372 79636
rect 140228 75744 140280 75750
rect 140228 75686 140280 75692
rect 140136 75676 140188 75682
rect 140136 75618 140188 75624
rect 140332 75562 140360 79630
rect 140424 76498 140452 79766
rect 140412 76492 140464 76498
rect 140412 76434 140464 76440
rect 140412 76356 140464 76362
rect 140412 76298 140464 76304
rect 140056 75534 140360 75562
rect 140056 68474 140084 75534
rect 140136 74520 140188 74526
rect 140136 74462 140188 74468
rect 140044 68468 140096 68474
rect 140044 68410 140096 68416
rect 140044 67584 140096 67590
rect 140044 67526 140096 67532
rect 139952 67108 140004 67114
rect 139952 67050 140004 67056
rect 139860 27260 139912 27266
rect 139860 27202 139912 27208
rect 139676 27192 139728 27198
rect 139676 27134 139728 27140
rect 139584 14340 139636 14346
rect 139584 14282 139636 14288
rect 139492 11552 139544 11558
rect 139492 11494 139544 11500
rect 139400 6860 139452 6866
rect 139400 6802 139452 6808
rect 140056 3890 140084 67526
rect 140148 4010 140176 74462
rect 140424 64874 140452 76298
rect 140516 73137 140544 79784
rect 140654 79744 140682 80036
rect 140608 79716 140682 79744
rect 140608 75857 140636 79716
rect 140746 79676 140774 80036
rect 140838 79898 140866 80036
rect 140930 79971 140958 80036
rect 140916 79962 140972 79971
rect 140826 79892 140878 79898
rect 140916 79897 140972 79906
rect 140826 79834 140878 79840
rect 141022 79778 141050 80036
rect 141114 79830 141142 80036
rect 140976 79750 141050 79778
rect 141102 79824 141154 79830
rect 141102 79766 141154 79772
rect 141206 79778 141234 80036
rect 141298 79937 141326 80036
rect 141284 79928 141340 79937
rect 141284 79863 141340 79872
rect 141390 79812 141418 80036
rect 141482 79966 141510 80036
rect 141574 79971 141602 80036
rect 141470 79960 141522 79966
rect 141470 79902 141522 79908
rect 141560 79962 141616 79971
rect 141666 79966 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141560 79897 141616 79906
rect 141654 79960 141706 79966
rect 141654 79902 141706 79908
rect 141746 79960 141798 79966
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141942 79937 141970 80036
rect 141838 79902 141890 79908
rect 141928 79928 141984 79937
rect 142034 79898 142062 80036
rect 142126 79971 142154 80036
rect 142112 79962 142168 79971
rect 142218 79966 142246 80036
rect 142310 79966 142338 80036
rect 141928 79863 141984 79872
rect 142022 79892 142074 79898
rect 142112 79897 142168 79906
rect 142206 79960 142258 79966
rect 142206 79902 142258 79908
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142022 79834 142074 79840
rect 141700 79824 141752 79830
rect 141390 79784 141556 79812
rect 141206 79750 141326 79778
rect 140700 79648 140774 79676
rect 140872 79688 140924 79694
rect 140594 75848 140650 75857
rect 140594 75783 140650 75792
rect 140700 75585 140728 79648
rect 140976 79665 141004 79750
rect 141298 79744 141326 79750
rect 141298 79716 141372 79744
rect 141148 79688 141200 79694
rect 140872 79630 140924 79636
rect 140962 79656 141018 79665
rect 140884 78849 140912 79630
rect 141148 79630 141200 79636
rect 140962 79591 141018 79600
rect 141056 79552 141108 79558
rect 141056 79494 141108 79500
rect 140964 79484 141016 79490
rect 140964 79426 141016 79432
rect 140870 78840 140926 78849
rect 140870 78775 140926 78784
rect 140872 78668 140924 78674
rect 140872 78610 140924 78616
rect 140780 76084 140832 76090
rect 140780 76026 140832 76032
rect 140686 75576 140742 75585
rect 140686 75511 140742 75520
rect 140502 73128 140558 73137
rect 140502 73063 140558 73072
rect 140332 64846 140452 64874
rect 140332 25974 140360 64846
rect 140320 25968 140372 25974
rect 140320 25910 140372 25916
rect 140136 4004 140188 4010
rect 140136 3946 140188 3952
rect 140792 3942 140820 76026
rect 140780 3936 140832 3942
rect 140056 3862 140176 3890
rect 140780 3878 140832 3884
rect 140884 3874 140912 78610
rect 140044 3596 140096 3602
rect 140044 3538 140096 3544
rect 139032 3324 139084 3330
rect 139032 3266 139084 3272
rect 140056 480 140084 3538
rect 140148 3466 140176 3862
rect 140872 3868 140924 3874
rect 140872 3810 140924 3816
rect 140976 3602 141004 79426
rect 141068 78402 141096 79494
rect 141056 78396 141108 78402
rect 141056 78338 141108 78344
rect 141056 78260 141108 78266
rect 141056 78202 141108 78208
rect 141068 5166 141096 78202
rect 141160 76090 141188 79630
rect 141240 79620 141292 79626
rect 141240 79562 141292 79568
rect 141148 76084 141200 76090
rect 141148 76026 141200 76032
rect 141148 75948 141200 75954
rect 141148 75890 141200 75896
rect 141160 28490 141188 75890
rect 141252 28558 141280 79562
rect 141344 28626 141372 79716
rect 141422 79656 141478 79665
rect 141422 79591 141478 79600
rect 141436 32910 141464 79591
rect 141528 78674 141556 79784
rect 141606 79792 141662 79801
rect 141700 79766 141752 79772
rect 141974 79792 142030 79801
rect 141606 79727 141662 79736
rect 141516 78668 141568 78674
rect 141516 78610 141568 78616
rect 141620 78266 141648 79727
rect 141608 78260 141660 78266
rect 141608 78202 141660 78208
rect 141606 78160 141662 78169
rect 141606 78095 141662 78104
rect 141620 70394 141648 78095
rect 141712 75954 141740 79766
rect 141884 79756 141936 79762
rect 141974 79727 142030 79736
rect 142068 79756 142120 79762
rect 141884 79698 141936 79704
rect 141792 79688 141844 79694
rect 141792 79630 141844 79636
rect 141804 76401 141832 79630
rect 141790 76392 141846 76401
rect 141790 76327 141846 76336
rect 141700 75948 141752 75954
rect 141700 75890 141752 75896
rect 141896 73982 141924 79698
rect 141988 77081 142016 79727
rect 142402 79744 142430 80036
rect 142494 79903 142522 80036
rect 142480 79894 142536 79903
rect 142480 79829 142536 79838
rect 142402 79716 142476 79744
rect 142068 79698 142120 79704
rect 142080 77926 142108 79698
rect 142342 79656 142398 79665
rect 142342 79591 142398 79600
rect 142068 77920 142120 77926
rect 142068 77862 142120 77868
rect 141974 77072 142030 77081
rect 141974 77007 142030 77016
rect 142252 74180 142304 74186
rect 142252 74122 142304 74128
rect 141884 73976 141936 73982
rect 141884 73918 141936 73924
rect 141528 70366 141648 70394
rect 141424 32904 141476 32910
rect 141424 32846 141476 32852
rect 141528 32842 141556 70366
rect 141516 32836 141568 32842
rect 141516 32778 141568 32784
rect 141332 28620 141384 28626
rect 141332 28562 141384 28568
rect 141240 28552 141292 28558
rect 141240 28494 141292 28500
rect 141148 28484 141200 28490
rect 141148 28426 141200 28432
rect 142264 7886 142292 74122
rect 142252 7880 142304 7886
rect 142252 7822 142304 7828
rect 141056 5160 141108 5166
rect 141056 5102 141108 5108
rect 142356 3913 142384 79591
rect 142448 17882 142476 79716
rect 142586 79608 142614 80036
rect 142678 79898 142706 80036
rect 142770 79898 142798 80036
rect 142666 79892 142718 79898
rect 142666 79834 142718 79840
rect 142758 79892 142810 79898
rect 142758 79834 142810 79840
rect 142862 79744 142890 80036
rect 142954 79971 142982 80036
rect 142940 79962 142996 79971
rect 142940 79897 142996 79906
rect 143046 79744 143074 80036
rect 142816 79716 142890 79744
rect 143000 79716 143074 79744
rect 143138 79744 143166 80036
rect 143230 79898 143258 80036
rect 143218 79892 143270 79898
rect 143218 79834 143270 79840
rect 143322 79801 143350 80036
rect 143414 79937 143442 80036
rect 143506 79966 143534 80036
rect 143494 79960 143546 79966
rect 143400 79928 143456 79937
rect 143494 79902 143546 79908
rect 143598 79898 143626 80036
rect 143400 79863 143456 79872
rect 143586 79892 143638 79898
rect 143586 79834 143638 79840
rect 143690 79830 143718 80036
rect 143782 79898 143810 80036
rect 143770 79892 143822 79898
rect 143770 79834 143822 79840
rect 143448 79824 143500 79830
rect 143308 79792 143364 79801
rect 143138 79716 143212 79744
rect 143448 79766 143500 79772
rect 143678 79824 143730 79830
rect 143874 79778 143902 80036
rect 143966 79830 143994 80036
rect 144058 79898 144086 80036
rect 144150 79971 144178 80036
rect 144136 79962 144192 79971
rect 144046 79892 144098 79898
rect 144136 79897 144192 79906
rect 144046 79834 144098 79840
rect 143678 79766 143730 79772
rect 143308 79727 143364 79736
rect 142540 79580 142614 79608
rect 142712 79620 142764 79626
rect 142540 27130 142568 79580
rect 142712 79562 142764 79568
rect 142620 79484 142672 79490
rect 142620 79426 142672 79432
rect 142632 29986 142660 79426
rect 142724 33862 142752 79562
rect 142816 74186 142844 79716
rect 142896 79620 142948 79626
rect 142896 79562 142948 79568
rect 142908 77761 142936 79562
rect 142894 77752 142950 77761
rect 142894 77687 142950 77696
rect 143000 75914 143028 79716
rect 143080 79416 143132 79422
rect 143080 79358 143132 79364
rect 142908 75886 143028 75914
rect 142804 74180 142856 74186
rect 142804 74122 142856 74128
rect 142908 70394 142936 75886
rect 142988 73568 143040 73574
rect 142988 73510 143040 73516
rect 142816 70366 142936 70394
rect 142816 63034 142844 70366
rect 142804 63028 142856 63034
rect 142804 62970 142856 62976
rect 142712 33856 142764 33862
rect 142712 33798 142764 33804
rect 142620 29980 142672 29986
rect 142620 29922 142672 29928
rect 142528 27124 142580 27130
rect 142528 27066 142580 27072
rect 142436 17876 142488 17882
rect 142436 17818 142488 17824
rect 142434 4040 142490 4049
rect 142434 3975 142490 3984
rect 142342 3904 142398 3913
rect 142342 3839 142398 3848
rect 140964 3596 141016 3602
rect 140964 3538 141016 3544
rect 140136 3460 140188 3466
rect 140136 3402 140188 3408
rect 141240 3188 141292 3194
rect 141240 3130 141292 3136
rect 141252 480 141280 3130
rect 142448 480 142476 3975
rect 143000 3398 143028 73510
rect 142988 3392 143040 3398
rect 142988 3334 143040 3340
rect 143092 3233 143120 79358
rect 143184 77178 143212 79716
rect 143264 79688 143316 79694
rect 143264 79630 143316 79636
rect 143172 77172 143224 77178
rect 143172 77114 143224 77120
rect 143276 76673 143304 79630
rect 143262 76664 143318 76673
rect 143262 76599 143318 76608
rect 143460 74089 143488 79766
rect 143828 79750 143902 79778
rect 143954 79824 144006 79830
rect 143954 79766 144006 79772
rect 144092 79756 144144 79762
rect 143540 79688 143592 79694
rect 143592 79648 143672 79676
rect 143828 79665 143856 79750
rect 144242 79744 144270 80036
rect 144334 79898 144362 80036
rect 144322 79892 144374 79898
rect 144322 79834 144374 79840
rect 144426 79778 144454 80036
rect 144518 79937 144546 80036
rect 144504 79928 144560 79937
rect 144504 79863 144560 79872
rect 144092 79698 144144 79704
rect 144196 79716 144270 79744
rect 144380 79750 144454 79778
rect 144610 79778 144638 80036
rect 144702 79971 144730 80036
rect 144688 79962 144744 79971
rect 144688 79897 144744 79906
rect 144794 79830 144822 80036
rect 144886 79966 144914 80036
rect 144978 79966 145006 80036
rect 145070 79966 145098 80036
rect 145162 79966 145190 80036
rect 145254 79966 145282 80036
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144966 79960 145018 79966
rect 144966 79902 145018 79908
rect 145058 79960 145110 79966
rect 145058 79902 145110 79908
rect 145150 79960 145202 79966
rect 145150 79902 145202 79908
rect 145242 79960 145294 79966
rect 145242 79902 145294 79908
rect 144782 79824 144834 79830
rect 144610 79750 144684 79778
rect 145346 79801 145374 80036
rect 145438 79830 145466 80036
rect 145530 79937 145558 80036
rect 145622 79966 145650 80036
rect 145714 79966 145742 80036
rect 145610 79960 145662 79966
rect 145516 79928 145572 79937
rect 145610 79902 145662 79908
rect 145702 79960 145754 79966
rect 145702 79902 145754 79908
rect 145516 79863 145572 79872
rect 145426 79824 145478 79830
rect 144782 79766 144834 79772
rect 145332 79792 145388 79801
rect 143908 79688 143960 79694
rect 143540 79630 143592 79636
rect 143540 79416 143592 79422
rect 143540 79358 143592 79364
rect 143552 79218 143580 79358
rect 143540 79212 143592 79218
rect 143540 79154 143592 79160
rect 143446 74080 143502 74089
rect 143446 74015 143502 74024
rect 143644 4146 143672 79648
rect 143814 79656 143870 79665
rect 143908 79630 143960 79636
rect 143814 79591 143870 79600
rect 143816 79484 143868 79490
rect 143816 79426 143868 79432
rect 143828 77217 143856 79426
rect 143814 77208 143870 77217
rect 143814 77143 143870 77152
rect 143724 76832 143776 76838
rect 143724 76774 143776 76780
rect 143736 6730 143764 76774
rect 143814 76664 143870 76673
rect 143814 76599 143870 76608
rect 143828 6798 143856 76599
rect 143920 12442 143948 79630
rect 144000 79552 144052 79558
rect 144000 79494 144052 79500
rect 143908 12436 143960 12442
rect 143908 12378 143960 12384
rect 144012 11694 144040 79494
rect 144104 16250 144132 79698
rect 144196 78198 144224 79716
rect 144276 79620 144328 79626
rect 144276 79562 144328 79568
rect 144184 78192 144236 78198
rect 144184 78134 144236 78140
rect 144184 75948 144236 75954
rect 144184 75890 144236 75896
rect 144196 18902 144224 75890
rect 144288 33794 144316 79562
rect 144380 76838 144408 79750
rect 144458 79656 144514 79665
rect 144458 79591 144514 79600
rect 144368 76832 144420 76838
rect 144368 76774 144420 76780
rect 144368 76696 144420 76702
rect 144368 76638 144420 76644
rect 144380 70394 144408 76638
rect 144472 71774 144500 79591
rect 144552 79552 144604 79558
rect 144552 79494 144604 79500
rect 144564 77897 144592 79494
rect 144550 77888 144606 77897
rect 144550 77823 144606 77832
rect 144656 73953 144684 79750
rect 144920 79756 144972 79762
rect 144920 79698 144972 79704
rect 145012 79756 145064 79762
rect 145064 79716 145144 79744
rect 145426 79766 145478 79772
rect 145656 79824 145708 79830
rect 145656 79766 145708 79772
rect 145332 79727 145388 79736
rect 145012 79698 145064 79704
rect 144736 79620 144788 79626
rect 144736 79562 144788 79568
rect 144828 79620 144880 79626
rect 144828 79562 144880 79568
rect 144748 75954 144776 79562
rect 144840 76906 144868 79562
rect 144932 77858 144960 79698
rect 145012 79552 145064 79558
rect 145012 79494 145064 79500
rect 144920 77852 144972 77858
rect 144920 77794 144972 77800
rect 144828 76900 144880 76906
rect 144828 76842 144880 76848
rect 145024 76090 145052 79494
rect 145116 76106 145144 79716
rect 145286 79656 145342 79665
rect 145286 79591 145342 79600
rect 145380 79620 145432 79626
rect 145012 76084 145064 76090
rect 145116 76078 145236 76106
rect 145012 76026 145064 76032
rect 145104 76016 145156 76022
rect 144918 75984 144974 75993
rect 144736 75948 144788 75954
rect 145104 75958 145156 75964
rect 144918 75919 144974 75928
rect 144736 75890 144788 75896
rect 144642 73944 144698 73953
rect 144642 73879 144698 73888
rect 144472 71746 144592 71774
rect 144380 70366 144500 70394
rect 144276 33788 144328 33794
rect 144276 33730 144328 33736
rect 144184 18896 144236 18902
rect 144184 18838 144236 18844
rect 144092 16244 144144 16250
rect 144092 16186 144144 16192
rect 144000 11688 144052 11694
rect 144000 11630 144052 11636
rect 143816 6792 143868 6798
rect 143816 6734 143868 6740
rect 143724 6724 143776 6730
rect 143724 6666 143776 6672
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 143632 4140 143684 4146
rect 143632 4082 143684 4088
rect 143078 3224 143134 3233
rect 143078 3159 143134 3168
rect 143552 480 143580 4082
rect 144472 3194 144500 70366
rect 144564 3505 144592 71746
rect 144932 6594 144960 75919
rect 145012 73772 145064 73778
rect 145012 73714 145064 73720
rect 144920 6588 144972 6594
rect 144920 6530 144972 6536
rect 145024 6526 145052 73714
rect 145116 6662 145144 75958
rect 145208 14414 145236 76078
rect 145300 15162 145328 79591
rect 145380 79562 145432 79568
rect 145472 79620 145524 79626
rect 145472 79562 145524 79568
rect 145392 76022 145420 79562
rect 145380 76016 145432 76022
rect 145380 75958 145432 75964
rect 145484 75914 145512 79562
rect 145668 77294 145696 79766
rect 145806 79744 145834 80036
rect 145898 79966 145926 80036
rect 145886 79960 145938 79966
rect 145886 79902 145938 79908
rect 145990 79898 146018 80036
rect 146082 79937 146110 80036
rect 146174 79966 146202 80036
rect 146162 79960 146214 79966
rect 146068 79928 146124 79937
rect 145978 79892 146030 79898
rect 146162 79902 146214 79908
rect 146068 79863 146124 79872
rect 145978 79834 146030 79840
rect 145932 79756 145984 79762
rect 145806 79716 145880 79744
rect 145746 79656 145802 79665
rect 145746 79591 145748 79600
rect 145800 79591 145802 79600
rect 145748 79562 145800 79568
rect 145392 75886 145512 75914
rect 145576 77266 145696 77294
rect 145288 15156 145340 15162
rect 145288 15098 145340 15104
rect 145392 15094 145420 75886
rect 145472 72956 145524 72962
rect 145472 72898 145524 72904
rect 145484 20670 145512 72898
rect 145472 20664 145524 20670
rect 145472 20606 145524 20612
rect 145576 19922 145604 77266
rect 145656 76016 145708 76022
rect 145656 75958 145708 75964
rect 145668 20534 145696 75958
rect 145852 73778 145880 79716
rect 146266 79744 146294 80036
rect 146358 79971 146386 80036
rect 146344 79962 146400 79971
rect 146450 79966 146478 80036
rect 146344 79897 146400 79906
rect 146438 79960 146490 79966
rect 146438 79902 146490 79908
rect 146542 79903 146570 80036
rect 146634 79966 146662 80036
rect 146726 79966 146754 80036
rect 146622 79960 146674 79966
rect 146528 79894 146584 79903
rect 146622 79902 146674 79908
rect 146714 79960 146766 79966
rect 146714 79902 146766 79908
rect 146528 79829 146584 79838
rect 146818 79812 146846 80036
rect 146910 79898 146938 80036
rect 146898 79892 146950 79898
rect 146898 79834 146950 79840
rect 146772 79784 146846 79812
rect 146772 79744 146800 79784
rect 145932 79698 145984 79704
rect 146220 79716 146294 79744
rect 146680 79716 146800 79744
rect 147002 79744 147030 80036
rect 147094 79898 147122 80036
rect 147186 79966 147214 80036
rect 147278 79966 147306 80036
rect 147370 79971 147398 80036
rect 147174 79960 147226 79966
rect 147174 79902 147226 79908
rect 147266 79960 147318 79966
rect 147266 79902 147318 79908
rect 147356 79962 147412 79971
rect 147462 79966 147490 80036
rect 147554 79971 147582 80036
rect 147082 79892 147134 79898
rect 147356 79897 147412 79906
rect 147450 79960 147502 79966
rect 147450 79902 147502 79908
rect 147540 79962 147596 79971
rect 147540 79897 147596 79906
rect 147646 79898 147674 80036
rect 147082 79834 147134 79840
rect 147634 79892 147686 79898
rect 147634 79834 147686 79840
rect 147312 79824 147364 79830
rect 147310 79792 147312 79801
rect 147364 79792 147366 79801
rect 147002 79716 147076 79744
rect 147310 79727 147366 79736
rect 147586 79792 147642 79801
rect 147738 79744 147766 80036
rect 147830 79971 147858 80036
rect 147816 79962 147872 79971
rect 147922 79966 147950 80036
rect 147816 79897 147872 79906
rect 147910 79960 147962 79966
rect 147910 79902 147962 79908
rect 147586 79727 147642 79736
rect 145840 73772 145892 73778
rect 145840 73714 145892 73720
rect 145944 72962 145972 79698
rect 146024 79688 146076 79694
rect 146024 79630 146076 79636
rect 146036 75857 146064 79630
rect 146022 75848 146078 75857
rect 146022 75783 146078 75792
rect 146220 74225 146248 79716
rect 146298 79656 146354 79665
rect 146298 79591 146354 79600
rect 146484 79620 146536 79626
rect 146206 74216 146262 74225
rect 146206 74151 146262 74160
rect 145932 72956 145984 72962
rect 145932 72898 145984 72904
rect 145656 20528 145708 20534
rect 145656 20470 145708 20476
rect 145564 19916 145616 19922
rect 145564 19858 145616 19864
rect 145380 15088 145432 15094
rect 145380 15030 145432 15036
rect 145196 14408 145248 14414
rect 145196 14350 145248 14356
rect 145104 6656 145156 6662
rect 145104 6598 145156 6604
rect 145012 6520 145064 6526
rect 145012 6462 145064 6468
rect 145932 5024 145984 5030
rect 145932 4966 145984 4972
rect 144736 3528 144788 3534
rect 144550 3496 144606 3505
rect 144736 3470 144788 3476
rect 144550 3431 144606 3440
rect 144460 3188 144512 3194
rect 144460 3130 144512 3136
rect 144748 480 144776 3470
rect 145944 480 145972 4966
rect 146312 3738 146340 79591
rect 146484 79562 146536 79568
rect 146392 79552 146444 79558
rect 146392 79494 146444 79500
rect 146404 6458 146432 79494
rect 146496 76090 146524 79562
rect 146680 76158 146708 79716
rect 146852 79688 146904 79694
rect 146852 79630 146904 79636
rect 146760 79620 146812 79626
rect 146760 79562 146812 79568
rect 146668 76152 146720 76158
rect 146668 76094 146720 76100
rect 146484 76084 146536 76090
rect 146484 76026 146536 76032
rect 146668 76016 146720 76022
rect 146668 75958 146720 75964
rect 146484 75948 146536 75954
rect 146484 75890 146536 75896
rect 146576 75948 146628 75954
rect 146576 75890 146628 75896
rect 146392 6452 146444 6458
rect 146392 6394 146444 6400
rect 146496 6390 146524 75890
rect 146588 9586 146616 75890
rect 146680 12374 146708 75958
rect 146772 14958 146800 79562
rect 146864 76226 146892 79630
rect 146944 79620 146996 79626
rect 146944 79562 146996 79568
rect 146852 76220 146904 76226
rect 146852 76162 146904 76168
rect 146852 76084 146904 76090
rect 146852 76026 146904 76032
rect 146864 15026 146892 76026
rect 146956 17678 146984 79562
rect 147048 76294 147076 79716
rect 147220 79688 147272 79694
rect 147126 79656 147182 79665
rect 147220 79630 147272 79636
rect 147496 79688 147548 79694
rect 147496 79630 147548 79636
rect 147126 79591 147182 79600
rect 147036 76288 147088 76294
rect 147036 76230 147088 76236
rect 147036 76152 147088 76158
rect 147036 76094 147088 76100
rect 147048 17746 147076 76094
rect 147140 70394 147168 79591
rect 147232 75954 147260 79630
rect 147310 76256 147366 76265
rect 147310 76191 147366 76200
rect 147220 75948 147272 75954
rect 147220 75890 147272 75896
rect 147324 73914 147352 76191
rect 147508 75993 147536 79630
rect 147600 77217 147628 79727
rect 147692 79716 147766 79744
rect 147862 79792 147918 79801
rect 147862 79727 147918 79736
rect 147692 78470 147720 79716
rect 147770 79656 147826 79665
rect 147770 79591 147826 79600
rect 147680 78464 147732 78470
rect 147680 78406 147732 78412
rect 147680 77580 147732 77586
rect 147680 77522 147732 77528
rect 147586 77208 147642 77217
rect 147586 77143 147642 77152
rect 147692 76566 147720 77522
rect 147680 76560 147732 76566
rect 147680 76502 147732 76508
rect 147680 76424 147732 76430
rect 147680 76366 147732 76372
rect 147494 75984 147550 75993
rect 147494 75919 147550 75928
rect 147312 73908 147364 73914
rect 147312 73850 147364 73856
rect 147140 70366 147444 70394
rect 147416 64874 147444 70366
rect 147140 64846 147444 64874
rect 147140 17814 147168 64846
rect 147128 17808 147180 17814
rect 147128 17750 147180 17756
rect 147036 17740 147088 17746
rect 147036 17682 147088 17688
rect 146944 17672 146996 17678
rect 146944 17614 146996 17620
rect 146852 15020 146904 15026
rect 146852 14962 146904 14968
rect 146760 14952 146812 14958
rect 146760 14894 146812 14900
rect 146668 12368 146720 12374
rect 146668 12310 146720 12316
rect 146576 9580 146628 9586
rect 146576 9522 146628 9528
rect 146484 6384 146536 6390
rect 146484 6326 146536 6332
rect 147692 5098 147720 76366
rect 147784 9382 147812 79591
rect 147876 76702 147904 79727
rect 148014 79608 148042 80036
rect 148106 79676 148134 80036
rect 148198 79830 148226 80036
rect 148290 79966 148318 80036
rect 148278 79960 148330 79966
rect 148382 79937 148410 80036
rect 148278 79902 148330 79908
rect 148368 79928 148424 79937
rect 148368 79863 148424 79872
rect 148186 79824 148238 79830
rect 148186 79766 148238 79772
rect 148324 79824 148376 79830
rect 148324 79766 148376 79772
rect 148232 79688 148284 79694
rect 148106 79648 148180 79676
rect 148014 79580 148088 79608
rect 147956 79484 148008 79490
rect 147956 79426 148008 79432
rect 147968 77160 147996 79426
rect 148060 77586 148088 79580
rect 148048 77580 148100 77586
rect 148048 77522 148100 77528
rect 147968 77132 148088 77160
rect 147956 77036 148008 77042
rect 147956 76978 148008 76984
rect 147864 76696 147916 76702
rect 147864 76638 147916 76644
rect 147864 76560 147916 76566
rect 147864 76502 147916 76508
rect 147876 9518 147904 76502
rect 147864 9512 147916 9518
rect 147864 9454 147916 9460
rect 147968 9450 147996 76978
rect 148060 76770 148088 77132
rect 148048 76764 148100 76770
rect 148048 76706 148100 76712
rect 148046 76664 148102 76673
rect 148046 76599 148102 76608
rect 148060 24546 148088 76599
rect 148152 25906 148180 79648
rect 148232 79630 148284 79636
rect 148244 76888 148272 79630
rect 148336 79608 148364 79766
rect 148474 79744 148502 80036
rect 148566 79971 148594 80036
rect 148552 79962 148608 79971
rect 148552 79897 148608 79906
rect 148658 79744 148686 80036
rect 148474 79716 148548 79744
rect 148336 79580 148456 79608
rect 148324 79484 148376 79490
rect 148324 79426 148376 79432
rect 148336 78946 148364 79426
rect 148324 78940 148376 78946
rect 148324 78882 148376 78888
rect 148428 77042 148456 79580
rect 148416 77036 148468 77042
rect 148416 76978 148468 76984
rect 148244 76860 148456 76888
rect 148324 76764 148376 76770
rect 148324 76706 148376 76712
rect 148232 76696 148284 76702
rect 148232 76638 148284 76644
rect 148244 32774 148272 76638
rect 148232 32768 148284 32774
rect 148232 32710 148284 32716
rect 148336 32706 148364 76706
rect 148428 35426 148456 76860
rect 148520 76430 148548 79716
rect 148612 79716 148686 79744
rect 148612 76838 148640 79716
rect 148750 79642 148778 80036
rect 148842 79971 148870 80036
rect 148828 79962 148884 79971
rect 148828 79897 148884 79906
rect 148934 79898 148962 80036
rect 148922 79892 148974 79898
rect 148922 79834 148974 79840
rect 149026 79801 149054 80036
rect 149012 79792 149068 79801
rect 149012 79727 149068 79736
rect 149118 79676 149146 80036
rect 149210 79966 149238 80036
rect 149198 79960 149250 79966
rect 149198 79902 149250 79908
rect 149302 79830 149330 80036
rect 149290 79824 149342 79830
rect 149290 79766 149342 79772
rect 149394 79744 149422 80036
rect 149486 79971 149514 80036
rect 149472 79962 149528 79971
rect 149472 79897 149528 79906
rect 149578 79744 149606 80036
rect 149670 79898 149698 80036
rect 149658 79892 149710 79898
rect 149658 79834 149710 79840
rect 149762 79778 149790 80036
rect 149854 79966 149882 80036
rect 149946 79966 149974 80036
rect 150038 79966 150066 80036
rect 150130 79966 150158 80036
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149934 79960 149986 79966
rect 149934 79902 149986 79908
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 150118 79960 150170 79966
rect 150118 79902 150170 79908
rect 150222 79801 150250 80036
rect 150314 79971 150342 80036
rect 150300 79962 150356 79971
rect 150300 79897 150356 79906
rect 149716 79750 149790 79778
rect 150208 79792 150264 79801
rect 149888 79756 149940 79762
rect 149394 79716 149468 79744
rect 149578 79716 149652 79744
rect 148966 79656 149022 79665
rect 148750 79614 148824 79642
rect 148692 79552 148744 79558
rect 148692 79494 148744 79500
rect 148600 76832 148652 76838
rect 148704 76809 148732 79494
rect 148600 76774 148652 76780
rect 148690 76800 148746 76809
rect 148690 76735 148746 76744
rect 148796 76673 148824 79614
rect 148966 79591 149022 79600
rect 149072 79648 149146 79676
rect 148782 76664 148838 76673
rect 148782 76599 148838 76608
rect 148508 76424 148560 76430
rect 148508 76366 148560 76372
rect 148980 74534 149008 79591
rect 149072 76650 149100 79648
rect 149244 79620 149296 79626
rect 149244 79562 149296 79568
rect 149152 79552 149204 79558
rect 149152 79494 149204 79500
rect 149164 76974 149192 79494
rect 149256 77042 149284 79562
rect 149336 79552 149388 79558
rect 149336 79494 149388 79500
rect 149244 77036 149296 77042
rect 149244 76978 149296 76984
rect 149152 76968 149204 76974
rect 149152 76910 149204 76916
rect 149244 76764 149296 76770
rect 149244 76706 149296 76712
rect 149072 76622 149192 76650
rect 148980 74506 149100 74534
rect 148416 35420 148468 35426
rect 148416 35362 148468 35368
rect 148324 32700 148376 32706
rect 148324 32642 148376 32648
rect 148140 25900 148192 25906
rect 148140 25842 148192 25848
rect 148048 24540 148100 24546
rect 148048 24482 148100 24488
rect 147956 9444 148008 9450
rect 147956 9386 148008 9392
rect 147772 9376 147824 9382
rect 147772 9318 147824 9324
rect 149072 7818 149100 74506
rect 149164 9314 149192 76622
rect 149152 9308 149204 9314
rect 149152 9250 149204 9256
rect 149256 9110 149284 76706
rect 149348 9178 149376 79494
rect 149440 9246 149468 79716
rect 149520 77308 149572 77314
rect 149520 77250 149572 77256
rect 149532 14890 149560 77250
rect 149624 77058 149652 79716
rect 149716 77314 149744 79750
rect 149888 79698 149940 79704
rect 149980 79756 150032 79762
rect 149980 79698 150032 79704
rect 150072 79756 150124 79762
rect 150208 79727 150264 79736
rect 150072 79698 150124 79704
rect 149796 79688 149848 79694
rect 149796 79630 149848 79636
rect 149704 77308 149756 77314
rect 149704 77250 149756 77256
rect 149624 77030 149744 77058
rect 149612 76968 149664 76974
rect 149612 76910 149664 76916
rect 149624 61470 149652 76910
rect 149716 72758 149744 77030
rect 149704 72752 149756 72758
rect 149704 72694 149756 72700
rect 149808 72690 149836 79630
rect 149900 76770 149928 79698
rect 149992 78169 150020 79698
rect 149978 78160 150034 78169
rect 149978 78095 150034 78104
rect 150084 77353 150112 79698
rect 150406 79676 150434 80036
rect 150498 79966 150526 80036
rect 150590 79966 150618 80036
rect 150486 79960 150538 79966
rect 150486 79902 150538 79908
rect 150578 79960 150630 79966
rect 150578 79902 150630 79908
rect 150682 79778 150710 80036
rect 150774 79966 150802 80036
rect 150762 79960 150814 79966
rect 150866 79937 150894 80036
rect 150958 79966 150986 80036
rect 150946 79960 150998 79966
rect 150762 79902 150814 79908
rect 150852 79928 150908 79937
rect 150946 79902 150998 79908
rect 151050 79898 151078 80036
rect 150852 79863 150908 79872
rect 151038 79892 151090 79898
rect 151038 79834 151090 79840
rect 150360 79648 150434 79676
rect 150636 79750 150710 79778
rect 150808 79824 150860 79830
rect 150808 79766 150860 79772
rect 150164 79620 150216 79626
rect 150164 79562 150216 79568
rect 150070 77344 150126 77353
rect 150070 77279 150126 77288
rect 149980 77036 150032 77042
rect 149980 76978 150032 76984
rect 149888 76764 149940 76770
rect 149888 76706 149940 76712
rect 149992 72826 150020 76978
rect 150176 76974 150204 79562
rect 150360 77382 150388 79648
rect 150440 79552 150492 79558
rect 150440 79494 150492 79500
rect 150452 78606 150480 79494
rect 150440 78600 150492 78606
rect 150440 78542 150492 78548
rect 150530 78160 150586 78169
rect 150530 78095 150586 78104
rect 150348 77376 150400 77382
rect 150348 77318 150400 77324
rect 150164 76968 150216 76974
rect 150164 76910 150216 76916
rect 150440 76016 150492 76022
rect 150440 75958 150492 75964
rect 149980 72820 150032 72826
rect 149980 72762 150032 72768
rect 149796 72684 149848 72690
rect 149796 72626 149848 72632
rect 149612 61464 149664 61470
rect 149612 61406 149664 61412
rect 149520 14884 149572 14890
rect 149520 14826 149572 14832
rect 149428 9240 149480 9246
rect 149428 9182 149480 9188
rect 149336 9172 149388 9178
rect 149336 9114 149388 9120
rect 149244 9104 149296 9110
rect 149244 9046 149296 9052
rect 149060 7812 149112 7818
rect 149060 7754 149112 7760
rect 150452 7750 150480 75958
rect 150544 10470 150572 78095
rect 150636 76022 150664 79750
rect 150716 79688 150768 79694
rect 150716 79630 150768 79636
rect 150624 76016 150676 76022
rect 150624 75958 150676 75964
rect 150624 75200 150676 75206
rect 150624 75142 150676 75148
rect 150636 12238 150664 75142
rect 150728 12306 150756 79630
rect 150820 75410 150848 79766
rect 150900 79756 150952 79762
rect 151142 79744 151170 80036
rect 150900 79698 150952 79704
rect 151096 79716 151170 79744
rect 150808 75404 150860 75410
rect 150808 75346 150860 75352
rect 150808 75268 150860 75274
rect 150808 75210 150860 75216
rect 150820 20602 150848 75210
rect 150912 32638 150940 79698
rect 150992 79620 151044 79626
rect 150992 79562 151044 79568
rect 151004 57322 151032 79562
rect 151096 75206 151124 79716
rect 151234 79642 151262 80036
rect 151326 79898 151354 80036
rect 151418 79966 151446 80036
rect 151510 79971 151538 80036
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151496 79962 151552 79971
rect 151314 79892 151366 79898
rect 151496 79897 151552 79906
rect 151314 79834 151366 79840
rect 151602 79812 151630 80036
rect 151358 79792 151414 79801
rect 151556 79784 151630 79812
rect 151694 79801 151722 80036
rect 151680 79792 151736 79801
rect 151358 79727 151414 79736
rect 151452 79756 151504 79762
rect 151188 79614 151262 79642
rect 151188 75274 151216 79614
rect 151268 79552 151320 79558
rect 151268 79494 151320 79500
rect 151176 75268 151228 75274
rect 151176 75210 151228 75216
rect 151084 75200 151136 75206
rect 151084 75142 151136 75148
rect 151280 70394 151308 79494
rect 151372 72622 151400 79727
rect 151452 79698 151504 79704
rect 151464 78742 151492 79698
rect 151452 78736 151504 78742
rect 151556 78713 151584 79784
rect 151680 79727 151736 79736
rect 151786 79676 151814 80036
rect 151878 79937 151906 80036
rect 151864 79928 151920 79937
rect 151864 79863 151920 79872
rect 151970 79812 151998 80036
rect 151740 79648 151814 79676
rect 151924 79784 151998 79812
rect 151740 78849 151768 79648
rect 151820 79552 151872 79558
rect 151820 79494 151872 79500
rect 151726 78840 151782 78849
rect 151726 78775 151782 78784
rect 151452 78678 151504 78684
rect 151542 78704 151598 78713
rect 151542 78639 151598 78648
rect 151360 72616 151412 72622
rect 151360 72558 151412 72564
rect 151096 70366 151308 70394
rect 151096 60246 151124 70366
rect 151084 60240 151136 60246
rect 151084 60182 151136 60188
rect 150992 57316 151044 57322
rect 150992 57258 151044 57264
rect 150900 32632 150952 32638
rect 150900 32574 150952 32580
rect 150808 20596 150860 20602
rect 150808 20538 150860 20544
rect 150716 12300 150768 12306
rect 150716 12242 150768 12248
rect 150624 12232 150676 12238
rect 150624 12174 150676 12180
rect 151832 12170 151860 79494
rect 151924 78946 151952 79784
rect 152062 79744 152090 80036
rect 152154 79966 152182 80036
rect 152142 79960 152194 79966
rect 152142 79902 152194 79908
rect 152246 79898 152274 80036
rect 152234 79892 152286 79898
rect 152234 79834 152286 79840
rect 152338 79744 152366 80036
rect 152430 79966 152458 80036
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152062 79716 152136 79744
rect 152004 79620 152056 79626
rect 152004 79562 152056 79568
rect 151912 78940 151964 78946
rect 151912 78882 151964 78888
rect 151910 78704 151966 78713
rect 151910 78639 151966 78648
rect 151924 75138 151952 78639
rect 151912 75132 151964 75138
rect 151912 75074 151964 75080
rect 151912 74996 151964 75002
rect 151912 74938 151964 74944
rect 151924 13462 151952 74938
rect 152016 16182 152044 79562
rect 152108 78810 152136 79716
rect 152200 79716 152366 79744
rect 152096 78804 152148 78810
rect 152096 78746 152148 78752
rect 152200 78010 152228 79716
rect 152522 79676 152550 80036
rect 152614 79937 152642 80036
rect 152600 79928 152656 79937
rect 152600 79863 152656 79872
rect 152706 79812 152734 80036
rect 152798 79830 152826 80036
rect 152890 79971 152918 80036
rect 152876 79962 152932 79971
rect 152876 79897 152932 79906
rect 152476 79648 152550 79676
rect 152660 79784 152734 79812
rect 152786 79824 152838 79830
rect 152280 79552 152332 79558
rect 152280 79494 152332 79500
rect 152108 77982 152228 78010
rect 152108 21690 152136 77982
rect 152188 77920 152240 77926
rect 152188 77862 152240 77868
rect 152200 77518 152228 77862
rect 152188 77512 152240 77518
rect 152188 77454 152240 77460
rect 152188 77308 152240 77314
rect 152292 77294 152320 79494
rect 152476 77314 152504 79648
rect 152556 79348 152608 79354
rect 152556 79290 152608 79296
rect 152568 78878 152596 79290
rect 152660 79082 152688 79784
rect 152982 79812 153010 80036
rect 152936 79801 153010 79812
rect 152786 79766 152838 79772
rect 152922 79792 153010 79801
rect 152978 79784 153010 79792
rect 153074 79744 153102 80036
rect 153166 79971 153194 80036
rect 153152 79962 153208 79971
rect 153258 79966 153286 80036
rect 153152 79897 153208 79906
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153200 79824 153252 79830
rect 153350 79778 153378 80036
rect 153442 79898 153470 80036
rect 153430 79892 153482 79898
rect 153430 79834 153482 79840
rect 153200 79766 153252 79772
rect 152922 79727 152978 79736
rect 153028 79716 153102 79744
rect 152740 79688 152792 79694
rect 153028 79642 153056 79716
rect 152740 79630 152792 79636
rect 152648 79076 152700 79082
rect 152648 79018 152700 79024
rect 152648 78940 152700 78946
rect 152648 78882 152700 78888
rect 152556 78872 152608 78878
rect 152556 78814 152608 78820
rect 152556 78192 152608 78198
rect 152556 78134 152608 78140
rect 152568 77858 152596 78134
rect 152556 77852 152608 77858
rect 152556 77794 152608 77800
rect 152464 77308 152516 77314
rect 152292 77266 152412 77294
rect 152188 77250 152240 77256
rect 152200 32570 152228 77250
rect 152280 76764 152332 76770
rect 152280 76706 152332 76712
rect 152188 32564 152240 32570
rect 152188 32506 152240 32512
rect 152292 32502 152320 76706
rect 152384 62966 152412 77266
rect 152464 77250 152516 77256
rect 152464 75132 152516 75138
rect 152464 75074 152516 75080
rect 152476 64530 152504 75074
rect 152660 70394 152688 78882
rect 152752 76770 152780 79630
rect 152936 79614 153056 79642
rect 153106 79656 153162 79665
rect 152832 77512 152884 77518
rect 152832 77454 152884 77460
rect 152740 76764 152792 76770
rect 152740 76706 152792 76712
rect 152568 70366 152688 70394
rect 152844 70394 152872 77454
rect 152936 77353 152964 79614
rect 153106 79591 153162 79600
rect 153120 79354 153148 79591
rect 153108 79348 153160 79354
rect 153108 79290 153160 79296
rect 153212 79218 153240 79766
rect 153304 79750 153378 79778
rect 153200 79212 153252 79218
rect 153200 79154 153252 79160
rect 153016 79076 153068 79082
rect 153016 79018 153068 79024
rect 152922 77344 152978 77353
rect 152922 77279 152978 77288
rect 153028 75002 153056 79018
rect 153200 78736 153252 78742
rect 153200 78678 153252 78684
rect 153108 77376 153160 77382
rect 153108 77318 153160 77324
rect 153120 75154 153148 77318
rect 153212 75274 153240 78678
rect 153200 75268 153252 75274
rect 153200 75210 153252 75216
rect 153120 75126 153240 75154
rect 153016 74996 153068 75002
rect 153016 74938 153068 74944
rect 153212 73846 153240 75126
rect 153200 73840 153252 73846
rect 153200 73782 153252 73788
rect 152844 70366 153056 70394
rect 152464 64524 152516 64530
rect 152464 64466 152516 64472
rect 152568 64462 152596 70366
rect 153028 64874 153056 70366
rect 152752 64846 153056 64874
rect 152556 64456 152608 64462
rect 152556 64398 152608 64404
rect 152372 62960 152424 62966
rect 152372 62902 152424 62908
rect 152464 61396 152516 61402
rect 152464 61338 152516 61344
rect 152280 32496 152332 32502
rect 152280 32438 152332 32444
rect 152096 21684 152148 21690
rect 152096 21626 152148 21632
rect 152004 16176 152056 16182
rect 152004 16118 152056 16124
rect 151912 13456 151964 13462
rect 151912 13398 151964 13404
rect 151820 12164 151872 12170
rect 151820 12106 151872 12112
rect 150532 10464 150584 10470
rect 150532 10406 150584 10412
rect 150440 7744 150492 7750
rect 150440 7686 150492 7692
rect 149520 6316 149572 6322
rect 149520 6258 149572 6264
rect 147680 5092 147732 5098
rect 147680 5034 147732 5040
rect 147036 4208 147088 4214
rect 147036 4150 147088 4156
rect 146944 4140 146996 4146
rect 146944 4082 146996 4088
rect 146850 4040 146906 4049
rect 146850 3975 146906 3984
rect 146300 3732 146352 3738
rect 146300 3674 146352 3680
rect 146864 3641 146892 3975
rect 146956 3806 146984 4082
rect 147048 3806 147076 4150
rect 146944 3800 146996 3806
rect 146944 3742 146996 3748
rect 147036 3800 147088 3806
rect 147036 3742 147088 3748
rect 146850 3632 146906 3641
rect 146850 3567 146906 3576
rect 147036 3392 147088 3398
rect 147220 3392 147272 3398
rect 147088 3340 147220 3346
rect 147036 3334 147272 3340
rect 147048 3318 147260 3334
rect 147128 3256 147180 3262
rect 147128 3198 147180 3204
rect 147140 480 147168 3198
rect 148324 3120 148376 3126
rect 148324 3062 148376 3068
rect 148336 480 148364 3062
rect 149532 480 149560 6258
rect 151820 4140 151872 4146
rect 151820 4082 151872 4088
rect 150624 4072 150676 4078
rect 150624 4014 150676 4020
rect 150636 480 150664 4014
rect 151832 480 151860 4082
rect 152476 4078 152504 61338
rect 152464 4072 152516 4078
rect 152464 4014 152516 4020
rect 152752 2990 152780 64846
rect 153304 13394 153332 79750
rect 153534 79744 153562 80036
rect 153488 79716 153562 79744
rect 153384 79688 153436 79694
rect 153384 79630 153436 79636
rect 153396 78674 153424 79630
rect 153384 78668 153436 78674
rect 153384 78610 153436 78616
rect 153384 77376 153436 77382
rect 153384 77318 153436 77324
rect 153292 13388 153344 13394
rect 153292 13330 153344 13336
rect 153396 13190 153424 77318
rect 153488 13326 153516 79716
rect 153626 79676 153654 80036
rect 153718 79966 153746 80036
rect 153706 79960 153758 79966
rect 153706 79902 153758 79908
rect 153810 79898 153838 80036
rect 153902 79966 153930 80036
rect 153890 79960 153942 79966
rect 153890 79902 153942 79908
rect 153798 79892 153850 79898
rect 153798 79834 153850 79840
rect 153994 79812 154022 80036
rect 153948 79801 154022 79812
rect 153934 79792 154022 79801
rect 153752 79756 153804 79762
rect 153752 79698 153804 79704
rect 153844 79756 153896 79762
rect 153990 79784 154022 79792
rect 153934 79727 153990 79736
rect 153844 79698 153896 79704
rect 153580 79648 153654 79676
rect 153580 16114 153608 79648
rect 153660 78668 153712 78674
rect 153660 78610 153712 78616
rect 153672 50454 153700 78610
rect 153764 60178 153792 79698
rect 153856 77294 153884 79698
rect 154086 79676 154114 80036
rect 154178 79898 154206 80036
rect 154270 79966 154298 80036
rect 154258 79960 154310 79966
rect 154258 79902 154310 79908
rect 154166 79892 154218 79898
rect 154166 79834 154218 79840
rect 154212 79756 154264 79762
rect 154362 79744 154390 80036
rect 154454 79812 154482 80036
rect 154546 79937 154574 80036
rect 154638 79966 154666 80036
rect 154626 79960 154678 79966
rect 154532 79928 154588 79937
rect 154626 79902 154678 79908
rect 154532 79863 154588 79872
rect 154454 79801 154528 79812
rect 154454 79792 154542 79801
rect 154454 79784 154486 79792
rect 154362 79716 154436 79744
rect 154730 79744 154758 80036
rect 154822 79778 154850 80036
rect 154914 79898 154942 80036
rect 154902 79892 154954 79898
rect 154902 79834 154954 79840
rect 154822 79750 154896 79778
rect 154486 79727 154542 79736
rect 154212 79698 154264 79704
rect 154086 79648 154160 79676
rect 154028 79552 154080 79558
rect 154028 79494 154080 79500
rect 154040 77450 154068 79494
rect 154028 77444 154080 77450
rect 154028 77386 154080 77392
rect 154132 77382 154160 79648
rect 154120 77376 154172 77382
rect 154120 77318 154172 77324
rect 154224 77314 154252 79698
rect 154408 79665 154436 79716
rect 154684 79716 154758 79744
rect 154488 79688 154540 79694
rect 154394 79656 154450 79665
rect 154488 79630 154540 79636
rect 154580 79688 154632 79694
rect 154580 79630 154632 79636
rect 154394 79591 154450 79600
rect 154396 78804 154448 78810
rect 154396 78746 154448 78752
rect 154212 77308 154264 77314
rect 153856 77266 153976 77294
rect 153948 77194 153976 77266
rect 154212 77250 154264 77256
rect 153948 77166 154252 77194
rect 154120 75268 154172 75274
rect 154120 75210 154172 75216
rect 153752 60172 153804 60178
rect 153752 60114 153804 60120
rect 153660 50448 153712 50454
rect 153660 50390 153712 50396
rect 154132 28422 154160 75210
rect 154224 70394 154252 77166
rect 154408 74534 154436 78746
rect 154500 77518 154528 79630
rect 154592 79082 154620 79630
rect 154580 79076 154632 79082
rect 154580 79018 154632 79024
rect 154684 77586 154712 79716
rect 154764 79620 154816 79626
rect 154764 79562 154816 79568
rect 154672 77580 154724 77586
rect 154672 77522 154724 77528
rect 154488 77512 154540 77518
rect 154488 77454 154540 77460
rect 154672 77444 154724 77450
rect 154672 77386 154724 77392
rect 154408 74506 154528 74534
rect 154500 72554 154528 74506
rect 154488 72548 154540 72554
rect 154488 72490 154540 72496
rect 154224 70366 154436 70394
rect 154120 28416 154172 28422
rect 154120 28358 154172 28364
rect 153568 16108 153620 16114
rect 153568 16050 153620 16056
rect 153476 13320 153528 13326
rect 153476 13262 153528 13268
rect 153384 13184 153436 13190
rect 153384 13126 153436 13132
rect 154212 6248 154264 6254
rect 154212 6190 154264 6196
rect 153016 3188 153068 3194
rect 153016 3130 153068 3136
rect 152740 2984 152792 2990
rect 152740 2926 152792 2932
rect 153028 480 153056 3130
rect 154224 480 154252 6190
rect 154408 5030 154436 70366
rect 154684 14686 154712 77386
rect 154776 14754 154804 79562
rect 154868 76702 154896 79750
rect 155006 79676 155034 80036
rect 155098 79744 155126 80036
rect 155190 79898 155218 80036
rect 155178 79892 155230 79898
rect 155178 79834 155230 79840
rect 155282 79744 155310 80036
rect 155374 79778 155402 80036
rect 155466 79898 155494 80036
rect 155454 79892 155506 79898
rect 155454 79834 155506 79840
rect 155374 79762 155448 79778
rect 155374 79756 155460 79762
rect 155374 79750 155408 79756
rect 155098 79716 155172 79744
rect 155006 79648 155080 79676
rect 154948 78804 155000 78810
rect 154948 78746 155000 78752
rect 154856 76696 154908 76702
rect 154856 76638 154908 76644
rect 154856 76560 154908 76566
rect 154856 76502 154908 76508
rect 154764 14748 154816 14754
rect 154764 14690 154816 14696
rect 154672 14680 154724 14686
rect 154672 14622 154724 14628
rect 154868 14618 154896 76502
rect 154960 14822 154988 78746
rect 155052 28354 155080 79648
rect 155144 78810 155172 79716
rect 155236 79716 155310 79744
rect 155132 78804 155184 78810
rect 155132 78746 155184 78752
rect 155236 78656 155264 79716
rect 155408 79698 155460 79704
rect 155558 79676 155586 80036
rect 155650 79744 155678 80036
rect 155742 79937 155770 80036
rect 155834 79966 155862 80036
rect 155926 79966 155954 80036
rect 156018 79966 156046 80036
rect 156110 79966 156138 80036
rect 156202 79971 156230 80036
rect 155822 79960 155874 79966
rect 155728 79928 155784 79937
rect 155822 79902 155874 79908
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 156006 79960 156058 79966
rect 156006 79902 156058 79908
rect 156098 79960 156150 79966
rect 156098 79902 156150 79908
rect 156188 79962 156244 79971
rect 156188 79897 156244 79906
rect 156294 79898 156322 80036
rect 156386 79971 156414 80036
rect 156372 79962 156428 79971
rect 156478 79966 156506 80036
rect 155728 79863 155784 79872
rect 156282 79892 156334 79898
rect 156372 79897 156428 79906
rect 156466 79960 156518 79966
rect 156466 79902 156518 79908
rect 156570 79898 156598 80036
rect 156662 79898 156690 80036
rect 156754 79966 156782 80036
rect 156742 79960 156794 79966
rect 156742 79902 156794 79908
rect 156282 79834 156334 79840
rect 156558 79892 156610 79898
rect 156558 79834 156610 79840
rect 156650 79892 156702 79898
rect 156650 79834 156702 79840
rect 156846 79778 156874 80036
rect 156938 79966 156966 80036
rect 157030 79966 157058 80036
rect 157122 79971 157150 80036
rect 156926 79960 156978 79966
rect 156926 79902 156978 79908
rect 157018 79960 157070 79966
rect 157018 79902 157070 79908
rect 157108 79962 157164 79971
rect 157214 79966 157242 80036
rect 157306 79971 157334 80036
rect 157108 79897 157164 79906
rect 157202 79960 157254 79966
rect 157202 79902 157254 79908
rect 157292 79962 157348 79971
rect 157292 79897 157348 79906
rect 157156 79824 157208 79830
rect 157076 79784 157156 79812
rect 157076 79778 157104 79784
rect 155776 79756 155828 79762
rect 155650 79716 155724 79744
rect 155558 79648 155632 79676
rect 155316 79620 155368 79626
rect 155316 79562 155368 79568
rect 155144 78628 155264 78656
rect 155144 71466 155172 78628
rect 155328 77450 155356 79562
rect 155500 79552 155552 79558
rect 155500 79494 155552 79500
rect 155512 77994 155540 79494
rect 155500 77988 155552 77994
rect 155500 77930 155552 77936
rect 155316 77444 155368 77450
rect 155316 77386 155368 77392
rect 155224 77376 155276 77382
rect 155224 77318 155276 77324
rect 155408 77376 155460 77382
rect 155408 77318 155460 77324
rect 155132 71460 155184 71466
rect 155132 71402 155184 71408
rect 155236 70394 155264 77318
rect 155420 76566 155448 77318
rect 155500 77308 155552 77314
rect 155500 77250 155552 77256
rect 155512 77092 155540 77250
rect 155604 77194 155632 79648
rect 155696 77382 155724 79716
rect 155776 79698 155828 79704
rect 155868 79756 155920 79762
rect 155868 79698 155920 79704
rect 156156 79750 156874 79778
rect 156984 79750 157104 79778
rect 157156 79766 157208 79772
rect 155684 77376 155736 77382
rect 155684 77318 155736 77324
rect 155788 77294 155816 79698
rect 155880 77654 155908 79698
rect 155958 79656 156014 79665
rect 155958 79591 156014 79600
rect 156052 79620 156104 79626
rect 155868 77648 155920 77654
rect 155868 77590 155920 77596
rect 155788 77266 155908 77294
rect 155604 77166 155816 77194
rect 155512 77064 155724 77092
rect 155408 76560 155460 76566
rect 155408 76502 155460 76508
rect 155236 70366 155632 70394
rect 155040 28348 155092 28354
rect 155040 28290 155092 28296
rect 154948 14816 155000 14822
rect 154948 14758 155000 14764
rect 154856 14612 154908 14618
rect 154856 14554 154908 14560
rect 155604 13258 155632 70366
rect 155696 65686 155724 77064
rect 155788 70394 155816 77166
rect 155880 76945 155908 77266
rect 155866 76936 155922 76945
rect 155866 76871 155922 76880
rect 155788 70366 155908 70394
rect 155684 65680 155736 65686
rect 155684 65622 155736 65628
rect 155592 13252 155644 13258
rect 155592 13194 155644 13200
rect 155880 7682 155908 70366
rect 155868 7676 155920 7682
rect 155868 7618 155920 7624
rect 155972 6322 156000 79591
rect 156052 79562 156104 79568
rect 156064 75070 156092 79562
rect 156052 75064 156104 75070
rect 156052 75006 156104 75012
rect 156052 74928 156104 74934
rect 156052 74870 156104 74876
rect 156064 12102 156092 74870
rect 156156 15910 156184 79750
rect 156328 79688 156380 79694
rect 156328 79630 156380 79636
rect 156420 79688 156472 79694
rect 156420 79630 156472 79636
rect 156512 79688 156564 79694
rect 156696 79688 156748 79694
rect 156512 79630 156564 79636
rect 156602 79656 156658 79665
rect 156236 79552 156288 79558
rect 156236 79494 156288 79500
rect 156248 75313 156276 79494
rect 156234 75304 156290 75313
rect 156234 75239 156290 75248
rect 156236 75200 156288 75206
rect 156236 75142 156288 75148
rect 156248 15978 156276 75142
rect 156340 16046 156368 79630
rect 156432 78810 156460 79630
rect 156420 78804 156472 78810
rect 156420 78746 156472 78752
rect 156420 77308 156472 77314
rect 156420 77250 156472 77256
rect 156432 26994 156460 77250
rect 156524 75206 156552 79630
rect 156696 79630 156748 79636
rect 156788 79688 156840 79694
rect 156984 79676 157012 79750
rect 156788 79630 156840 79636
rect 156938 79648 157012 79676
rect 156602 79591 156658 79600
rect 156512 75200 156564 75206
rect 156512 75142 156564 75148
rect 156512 75064 156564 75070
rect 156512 75006 156564 75012
rect 156524 29918 156552 75006
rect 156616 60110 156644 79591
rect 156708 77314 156736 79630
rect 156696 77308 156748 77314
rect 156696 77250 156748 77256
rect 156694 75168 156750 75177
rect 156694 75103 156750 75112
rect 156708 70394 156736 75103
rect 156800 74934 156828 79630
rect 156938 79540 156966 79648
rect 157064 79620 157116 79626
rect 157064 79562 157116 79568
rect 156938 79512 157012 79540
rect 156984 78713 157012 79512
rect 156970 78704 157026 78713
rect 156970 78639 157026 78648
rect 156972 78600 157024 78606
rect 156972 78542 157024 78548
rect 156788 74928 156840 74934
rect 156788 74870 156840 74876
rect 156708 70366 156828 70394
rect 156800 64874 156828 70366
rect 156984 68338 157012 78542
rect 157076 78062 157104 79562
rect 157156 79552 157208 79558
rect 157156 79494 157208 79500
rect 157248 79552 157300 79558
rect 157248 79494 157300 79500
rect 157064 78056 157116 78062
rect 157064 77998 157116 78004
rect 157168 75449 157196 79494
rect 157260 77296 157288 79494
rect 157398 79472 157426 80036
rect 157490 79898 157518 80036
rect 157478 79892 157530 79898
rect 157478 79834 157530 79840
rect 157582 79801 157610 80036
rect 157674 79898 157702 80036
rect 157766 79966 157794 80036
rect 157754 79960 157806 79966
rect 157754 79902 157806 79908
rect 157858 79898 157886 80036
rect 157662 79892 157714 79898
rect 157662 79834 157714 79840
rect 157846 79892 157898 79898
rect 157846 79834 157898 79840
rect 157568 79792 157624 79801
rect 157568 79727 157624 79736
rect 157798 79792 157854 79801
rect 157798 79727 157854 79736
rect 157950 79744 157978 80036
rect 158042 79812 158070 80036
rect 158134 79937 158162 80036
rect 158120 79928 158176 79937
rect 158120 79863 158176 79872
rect 158226 79830 158254 80036
rect 158318 79937 158346 80036
rect 158410 79966 158438 80036
rect 158398 79960 158450 79966
rect 158304 79928 158360 79937
rect 158398 79902 158450 79908
rect 158502 79898 158530 80036
rect 158594 79971 158622 80036
rect 158580 79962 158636 79971
rect 158686 79966 158714 80036
rect 158778 79966 158806 80036
rect 158304 79863 158360 79872
rect 158490 79892 158542 79898
rect 158580 79897 158636 79906
rect 158674 79960 158726 79966
rect 158674 79902 158726 79908
rect 158766 79960 158818 79966
rect 158766 79902 158818 79908
rect 158870 79898 158898 80036
rect 158962 79903 158990 80036
rect 158490 79834 158542 79840
rect 158858 79892 158910 79898
rect 158858 79834 158910 79840
rect 158948 79894 159004 79903
rect 159054 79898 159082 80036
rect 159146 79966 159174 80036
rect 159134 79960 159186 79966
rect 159134 79902 159186 79908
rect 159238 79898 159266 80036
rect 159330 79937 159358 80036
rect 159316 79928 159372 79937
rect 158214 79824 158266 79830
rect 158948 79829 159004 79838
rect 159042 79892 159094 79898
rect 159042 79834 159094 79840
rect 159226 79892 159278 79898
rect 159422 79898 159450 80036
rect 159514 79937 159542 80036
rect 159500 79928 159556 79937
rect 159316 79863 159372 79872
rect 159410 79892 159462 79898
rect 159226 79834 159278 79840
rect 159606 79898 159634 80036
rect 159500 79863 159556 79872
rect 159594 79892 159646 79898
rect 159410 79834 159462 79840
rect 159594 79834 159646 79840
rect 158042 79784 158116 79812
rect 157616 79620 157668 79626
rect 157616 79562 157668 79568
rect 157524 79552 157576 79558
rect 157524 79494 157576 79500
rect 157398 79444 157472 79472
rect 157444 77450 157472 79444
rect 157432 77444 157484 77450
rect 157432 77386 157484 77392
rect 157260 77268 157472 77296
rect 157340 75676 157392 75682
rect 157340 75618 157392 75624
rect 157154 75440 157210 75449
rect 157154 75375 157210 75384
rect 156972 68332 157024 68338
rect 156972 68274 157024 68280
rect 156708 64846 156828 64874
rect 156708 64394 156736 64846
rect 156696 64388 156748 64394
rect 156696 64330 156748 64336
rect 156604 60104 156656 60110
rect 156604 60046 156656 60052
rect 156512 29912 156564 29918
rect 156512 29854 156564 29860
rect 156420 26988 156472 26994
rect 156420 26930 156472 26936
rect 157352 17542 157380 75618
rect 157444 25838 157472 77268
rect 157536 29850 157564 79494
rect 157628 76770 157656 79562
rect 157708 79552 157760 79558
rect 157708 79494 157760 79500
rect 157720 79218 157748 79494
rect 157708 79212 157760 79218
rect 157708 79154 157760 79160
rect 157812 78946 157840 79727
rect 157950 79716 158024 79744
rect 157890 79656 157946 79665
rect 157890 79591 157892 79600
rect 157944 79591 157946 79600
rect 157892 79562 157944 79568
rect 157800 78940 157852 78946
rect 157800 78882 157852 78888
rect 157996 77602 158024 79716
rect 157720 77574 158024 77602
rect 157616 76764 157668 76770
rect 157616 76706 157668 76712
rect 157616 76628 157668 76634
rect 157616 76570 157668 76576
rect 157524 29844 157576 29850
rect 157524 29786 157576 29792
rect 157628 29782 157656 76570
rect 157720 57254 157748 77574
rect 157984 77444 158036 77450
rect 157984 77386 158036 77392
rect 157798 77344 157854 77353
rect 157798 77279 157854 77288
rect 157812 61402 157840 77279
rect 157892 76764 157944 76770
rect 157892 76706 157944 76712
rect 157904 67046 157932 76706
rect 157996 71398 158024 77386
rect 158088 76634 158116 79784
rect 158214 79766 158266 79772
rect 158444 79756 158496 79762
rect 158444 79698 158496 79704
rect 158812 79756 158864 79762
rect 159364 79756 159416 79762
rect 158864 79716 158944 79744
rect 158812 79698 158864 79704
rect 158168 79688 158220 79694
rect 158168 79630 158220 79636
rect 158076 76628 158128 76634
rect 158076 76570 158128 76576
rect 158180 75682 158208 79630
rect 158352 79620 158404 79626
rect 158352 79562 158404 79568
rect 158260 77580 158312 77586
rect 158260 77522 158312 77528
rect 158168 75676 158220 75682
rect 158168 75618 158220 75624
rect 157984 71392 158036 71398
rect 157984 71334 158036 71340
rect 158272 70394 158300 77522
rect 158364 74497 158392 79562
rect 158456 76673 158484 79698
rect 158718 79656 158774 79665
rect 158718 79591 158774 79600
rect 158628 77512 158680 77518
rect 158628 77454 158680 77460
rect 158442 76664 158498 76673
rect 158442 76599 158498 76608
rect 158350 74488 158406 74497
rect 158350 74423 158406 74432
rect 158640 72486 158668 77454
rect 158628 72480 158680 72486
rect 158628 72422 158680 72428
rect 158272 70366 158392 70394
rect 157892 67040 157944 67046
rect 157892 66982 157944 66988
rect 157800 61396 157852 61402
rect 157800 61338 157852 61344
rect 158364 58750 158392 70366
rect 158352 58744 158404 58750
rect 158352 58686 158404 58692
rect 157708 57248 157760 57254
rect 157708 57190 157760 57196
rect 157616 29776 157668 29782
rect 157616 29718 157668 29724
rect 157432 25832 157484 25838
rect 157432 25774 157484 25780
rect 157340 17536 157392 17542
rect 157340 17478 157392 17484
rect 156328 16040 156380 16046
rect 156328 15982 156380 15988
rect 156236 15972 156288 15978
rect 156236 15914 156288 15920
rect 156144 15904 156196 15910
rect 156144 15846 156196 15852
rect 156052 12096 156104 12102
rect 156052 12038 156104 12044
rect 158732 7614 158760 79591
rect 158916 77722 158944 79716
rect 159364 79698 159416 79704
rect 159548 79756 159600 79762
rect 159548 79698 159600 79704
rect 159088 79688 159140 79694
rect 159088 79630 159140 79636
rect 159180 79688 159232 79694
rect 159180 79630 159232 79636
rect 159270 79656 159326 79665
rect 158996 79620 159048 79626
rect 158996 79562 159048 79568
rect 158904 77716 158956 77722
rect 158904 77658 158956 77664
rect 158904 75948 158956 75954
rect 158904 75890 158956 75896
rect 158812 74996 158864 75002
rect 158812 74938 158864 74944
rect 158824 18766 158852 74938
rect 158916 21554 158944 75890
rect 159008 29714 159036 79562
rect 159100 75970 159128 79630
rect 159192 79014 159220 79630
rect 159270 79591 159326 79600
rect 159180 79008 159232 79014
rect 159180 78950 159232 78956
rect 159178 77888 159234 77897
rect 159178 77823 159234 77832
rect 159192 77790 159220 77823
rect 159180 77784 159232 77790
rect 159180 77726 159232 77732
rect 159100 75942 159220 75970
rect 159088 75744 159140 75750
rect 159088 75686 159140 75692
rect 159100 58682 159128 75686
rect 159192 60042 159220 75942
rect 159284 75002 159312 79591
rect 159376 78198 159404 79698
rect 159454 79656 159510 79665
rect 159454 79591 159510 79600
rect 159364 78192 159416 78198
rect 159364 78134 159416 78140
rect 159468 75954 159496 79591
rect 159456 75948 159508 75954
rect 159456 75890 159508 75896
rect 159272 74996 159324 75002
rect 159272 74938 159324 74944
rect 159560 70394 159588 79698
rect 159698 79676 159726 80036
rect 159790 79971 159818 80036
rect 159776 79962 159832 79971
rect 159882 79966 159910 80036
rect 159974 79966 160002 80036
rect 159776 79897 159832 79906
rect 159870 79960 159922 79966
rect 159870 79902 159922 79908
rect 159962 79960 160014 79966
rect 159962 79902 160014 79908
rect 160066 79898 160094 80036
rect 160158 79966 160186 80036
rect 160146 79960 160198 79966
rect 160250 79937 160278 80036
rect 160146 79902 160198 79908
rect 160236 79928 160292 79937
rect 160054 79892 160106 79898
rect 160236 79863 160292 79872
rect 160054 79834 160106 79840
rect 160342 79812 160370 80036
rect 159822 79792 159878 79801
rect 160158 79784 160370 79812
rect 160158 79778 160186 79784
rect 159822 79727 159878 79736
rect 160112 79750 160186 79778
rect 159698 79648 159772 79676
rect 159640 79552 159692 79558
rect 159640 79494 159692 79500
rect 159652 78606 159680 79494
rect 159640 78600 159692 78606
rect 159640 78542 159692 78548
rect 159640 77988 159692 77994
rect 159640 77930 159692 77936
rect 159284 70366 159588 70394
rect 159652 70394 159680 77930
rect 159744 75478 159772 79648
rect 159836 79642 159864 79727
rect 160112 79665 160140 79750
rect 160434 79744 160462 80036
rect 160526 79966 160554 80036
rect 160618 79966 160646 80036
rect 160514 79960 160566 79966
rect 160514 79902 160566 79908
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160710 79830 160738 80036
rect 160698 79824 160750 79830
rect 160698 79766 160750 79772
rect 160434 79716 160508 79744
rect 160098 79656 160154 79665
rect 159836 79614 159956 79642
rect 159824 79552 159876 79558
rect 159824 79494 159876 79500
rect 159836 75750 159864 79494
rect 159928 77586 159956 79614
rect 160008 79620 160060 79626
rect 160098 79591 160154 79600
rect 160192 79620 160244 79626
rect 160008 79562 160060 79568
rect 160192 79562 160244 79568
rect 159916 77580 159968 77586
rect 159916 77522 159968 77528
rect 159824 75744 159876 75750
rect 159824 75686 159876 75692
rect 159732 75472 159784 75478
rect 159732 75414 159784 75420
rect 159652 70366 159772 70394
rect 159284 68406 159312 70366
rect 159272 68400 159324 68406
rect 159272 68342 159324 68348
rect 159180 60036 159232 60042
rect 159180 59978 159232 59984
rect 159088 58676 159140 58682
rect 159088 58618 159140 58624
rect 159744 35358 159772 70366
rect 159732 35352 159784 35358
rect 159732 35294 159784 35300
rect 158996 29708 159048 29714
rect 158996 29650 159048 29656
rect 158904 21548 158956 21554
rect 158904 21490 158956 21496
rect 158812 18760 158864 18766
rect 158812 18702 158864 18708
rect 160020 17474 160048 79562
rect 160100 79552 160152 79558
rect 160100 79494 160152 79500
rect 160112 76634 160140 79494
rect 160100 76628 160152 76634
rect 160100 76570 160152 76576
rect 160100 76220 160152 76226
rect 160100 76162 160152 76168
rect 160112 75834 160140 76162
rect 160204 75993 160232 79562
rect 160376 79552 160428 79558
rect 160376 79494 160428 79500
rect 160388 79218 160416 79494
rect 160376 79212 160428 79218
rect 160376 79154 160428 79160
rect 160282 78840 160338 78849
rect 160282 78775 160338 78784
rect 160376 78804 160428 78810
rect 160190 75984 160246 75993
rect 160190 75919 160246 75928
rect 160112 75806 160232 75834
rect 160100 75744 160152 75750
rect 160100 75686 160152 75692
rect 160112 20194 160140 75686
rect 160204 20262 160232 75806
rect 160296 20398 160324 78775
rect 160376 78746 160428 78752
rect 160388 78470 160416 78746
rect 160376 78464 160428 78470
rect 160376 78406 160428 78412
rect 160374 75984 160430 75993
rect 160374 75919 160430 75928
rect 160284 20392 160336 20398
rect 160284 20334 160336 20340
rect 160192 20256 160244 20262
rect 160192 20198 160244 20204
rect 160100 20188 160152 20194
rect 160100 20130 160152 20136
rect 160388 20058 160416 75919
rect 160480 20330 160508 79716
rect 160802 79676 160830 80036
rect 160894 79937 160922 80036
rect 160986 79966 161014 80036
rect 160974 79960 161026 79966
rect 160880 79928 160936 79937
rect 161078 79937 161106 80036
rect 160974 79902 161026 79908
rect 161064 79928 161120 79937
rect 160880 79863 160936 79872
rect 161170 79898 161198 80036
rect 161262 79966 161290 80036
rect 161250 79960 161302 79966
rect 161250 79902 161302 79908
rect 161064 79863 161120 79872
rect 161158 79892 161210 79898
rect 161158 79834 161210 79840
rect 161354 79830 161382 80036
rect 161446 79971 161474 80036
rect 161432 79962 161488 79971
rect 161538 79966 161566 80036
rect 161432 79897 161488 79906
rect 161526 79960 161578 79966
rect 161630 79937 161658 80036
rect 161526 79902 161578 79908
rect 161616 79928 161672 79937
rect 161616 79863 161672 79872
rect 160928 79824 160980 79830
rect 160926 79792 160928 79801
rect 161342 79824 161394 79830
rect 160980 79792 160982 79801
rect 161342 79766 161394 79772
rect 160926 79727 160982 79736
rect 161572 79756 161624 79762
rect 161722 79744 161750 80036
rect 161814 79966 161842 80036
rect 161802 79960 161854 79966
rect 161802 79902 161854 79908
rect 161906 79744 161934 80036
rect 161572 79698 161624 79704
rect 161676 79716 161750 79744
rect 161860 79716 161934 79744
rect 160756 79648 160830 79676
rect 160928 79688 160980 79694
rect 160756 79472 160784 79648
rect 161112 79688 161164 79694
rect 160928 79630 160980 79636
rect 161110 79656 161112 79665
rect 161388 79688 161440 79694
rect 161164 79656 161166 79665
rect 160664 79444 160784 79472
rect 160560 79212 160612 79218
rect 160560 79154 160612 79160
rect 160572 76226 160600 79154
rect 160560 76220 160612 76226
rect 160560 76162 160612 76168
rect 160664 76158 160692 79444
rect 160744 79348 160796 79354
rect 160744 79290 160796 79296
rect 160756 79218 160784 79290
rect 160744 79212 160796 79218
rect 160744 79154 160796 79160
rect 160742 78704 160798 78713
rect 160940 78674 160968 79630
rect 161020 79620 161072 79626
rect 161388 79630 161440 79636
rect 161110 79591 161166 79600
rect 161296 79620 161348 79626
rect 161020 79562 161072 79568
rect 161296 79562 161348 79568
rect 160742 78639 160798 78648
rect 160928 78668 160980 78674
rect 160652 76152 160704 76158
rect 160652 76094 160704 76100
rect 160560 75948 160612 75954
rect 160560 75890 160612 75896
rect 160468 20324 160520 20330
rect 160468 20266 160520 20272
rect 160572 20126 160600 75890
rect 160650 75848 160706 75857
rect 160650 75783 160706 75792
rect 160664 28286 160692 75783
rect 160756 35222 160784 78639
rect 160928 78610 160980 78616
rect 160928 78124 160980 78130
rect 160928 78066 160980 78072
rect 160940 70394 160968 78066
rect 161032 75750 161060 79562
rect 161308 78169 161336 79562
rect 161294 78160 161350 78169
rect 161294 78095 161350 78104
rect 161400 76809 161428 79630
rect 161584 78810 161612 79698
rect 161572 78804 161624 78810
rect 161572 78746 161624 78752
rect 161572 78260 161624 78266
rect 161572 78202 161624 78208
rect 161386 76800 161442 76809
rect 161386 76735 161442 76744
rect 161480 75948 161532 75954
rect 161480 75890 161532 75896
rect 161020 75744 161072 75750
rect 161020 75686 161072 75692
rect 160940 70366 161152 70394
rect 160744 35216 160796 35222
rect 160744 35158 160796 35164
rect 160652 28280 160704 28286
rect 160652 28222 160704 28228
rect 160560 20120 160612 20126
rect 160560 20062 160612 20068
rect 160376 20052 160428 20058
rect 160376 19994 160428 20000
rect 160008 17468 160060 17474
rect 160008 17410 160060 17416
rect 158720 7608 158772 7614
rect 158720 7550 158772 7556
rect 155960 6316 156012 6322
rect 155960 6258 156012 6264
rect 160098 6216 160154 6225
rect 157800 6180 157852 6186
rect 160098 6151 160154 6160
rect 157800 6122 157852 6128
rect 154396 5024 154448 5030
rect 154396 4966 154448 4972
rect 155408 3392 155460 3398
rect 155408 3334 155460 3340
rect 155420 480 155448 3334
rect 156604 2984 156656 2990
rect 156604 2926 156656 2932
rect 156616 480 156644 2926
rect 157812 480 157840 6122
rect 158902 4856 158958 4865
rect 158902 4791 158958 4800
rect 158916 480 158944 4791
rect 160112 480 160140 6151
rect 161124 4146 161152 70366
rect 161492 6254 161520 75890
rect 161584 10402 161612 78202
rect 161676 78130 161704 79716
rect 161860 79642 161888 79716
rect 161998 79676 162026 80036
rect 162090 79830 162118 80036
rect 162182 79830 162210 80036
rect 162274 79966 162302 80036
rect 162262 79960 162314 79966
rect 162262 79902 162314 79908
rect 162366 79830 162394 80036
rect 162458 79966 162486 80036
rect 162550 79966 162578 80036
rect 162446 79960 162498 79966
rect 162446 79902 162498 79908
rect 162538 79960 162590 79966
rect 162538 79902 162590 79908
rect 162078 79824 162130 79830
rect 162078 79766 162130 79772
rect 162170 79824 162222 79830
rect 162170 79766 162222 79772
rect 162354 79824 162406 79830
rect 162354 79766 162406 79772
rect 162444 79826 162500 79835
rect 162642 79830 162670 80036
rect 162444 79761 162500 79770
rect 162630 79824 162682 79830
rect 162630 79766 162682 79772
rect 162734 79778 162762 80036
rect 162826 79966 162854 80036
rect 162814 79960 162866 79966
rect 162814 79902 162866 79908
rect 162918 79812 162946 80036
rect 162872 79801 162946 79812
rect 162858 79792 162946 79801
rect 162734 79750 162808 79778
rect 162124 79688 162176 79694
rect 161998 79648 162072 79676
rect 161860 79614 161934 79642
rect 161906 79540 161934 79614
rect 161860 79512 161934 79540
rect 161756 79484 161808 79490
rect 161756 79426 161808 79432
rect 161664 78124 161716 78130
rect 161664 78066 161716 78072
rect 161768 76158 161796 79426
rect 161756 76152 161808 76158
rect 161756 76094 161808 76100
rect 161756 76016 161808 76022
rect 161756 75958 161808 75964
rect 161664 73500 161716 73506
rect 161664 73442 161716 73448
rect 161676 12034 161704 73442
rect 161768 23050 161796 75958
rect 161860 32434 161888 79512
rect 161940 76152 161992 76158
rect 161940 76094 161992 76100
rect 161952 62898 161980 76094
rect 162044 76022 162072 79648
rect 162124 79630 162176 79636
rect 162216 79688 162268 79694
rect 162216 79630 162268 79636
rect 162308 79688 162360 79694
rect 162676 79688 162728 79694
rect 162308 79630 162360 79636
rect 162674 79656 162676 79665
rect 162728 79656 162730 79665
rect 162136 78266 162164 79630
rect 162124 78260 162176 78266
rect 162124 78202 162176 78208
rect 162124 77852 162176 77858
rect 162124 77794 162176 77800
rect 162032 76016 162084 76022
rect 162032 75958 162084 75964
rect 162030 75848 162086 75857
rect 162030 75783 162086 75792
rect 162044 64326 162072 75783
rect 162136 70394 162164 77794
rect 162228 75954 162256 79630
rect 162216 75948 162268 75954
rect 162216 75890 162268 75896
rect 162320 73506 162348 79630
rect 162492 79620 162544 79626
rect 162674 79591 162730 79600
rect 162492 79562 162544 79568
rect 162400 78668 162452 78674
rect 162400 78610 162452 78616
rect 162412 78266 162440 78610
rect 162400 78260 162452 78266
rect 162400 78202 162452 78208
rect 162504 77738 162532 79562
rect 162584 79552 162636 79558
rect 162584 79494 162636 79500
rect 162412 77710 162532 77738
rect 162412 75857 162440 77710
rect 162492 77648 162544 77654
rect 162492 77590 162544 77596
rect 162398 75848 162454 75857
rect 162398 75783 162454 75792
rect 162308 73500 162360 73506
rect 162308 73442 162360 73448
rect 162136 70366 162440 70394
rect 162032 64320 162084 64326
rect 162032 64262 162084 64268
rect 161940 62892 161992 62898
rect 161940 62834 161992 62840
rect 161848 32428 161900 32434
rect 161848 32370 161900 32376
rect 161756 23044 161808 23050
rect 161756 22986 161808 22992
rect 161664 12028 161716 12034
rect 161664 11970 161716 11976
rect 162412 11626 162440 70366
rect 162504 35290 162532 77590
rect 162596 75546 162624 79494
rect 162676 79484 162728 79490
rect 162676 79426 162728 79432
rect 162688 77897 162716 79426
rect 162674 77888 162730 77897
rect 162674 77823 162730 77832
rect 162780 75993 162808 79750
rect 162914 79784 162946 79792
rect 163010 79778 163038 80036
rect 163102 79966 163130 80036
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 163010 79750 163084 79778
rect 162858 79727 162914 79736
rect 162952 79688 163004 79694
rect 162872 79648 162952 79676
rect 162872 76265 162900 79648
rect 162952 79630 163004 79636
rect 162952 79552 163004 79558
rect 162952 79494 163004 79500
rect 162964 78305 162992 79494
rect 162950 78296 163006 78305
rect 162950 78231 163006 78240
rect 162952 78192 163004 78198
rect 162952 78134 163004 78140
rect 162964 77994 162992 78134
rect 162952 77988 163004 77994
rect 162952 77930 163004 77936
rect 162858 76256 162914 76265
rect 162858 76191 162914 76200
rect 162860 76084 162912 76090
rect 162860 76026 162912 76032
rect 162952 76084 163004 76090
rect 162952 76026 163004 76032
rect 162766 75984 162822 75993
rect 162766 75919 162822 75928
rect 162584 75540 162636 75546
rect 162584 75482 162636 75488
rect 162492 35284 162544 35290
rect 162492 35226 162544 35232
rect 162872 13122 162900 76026
rect 162964 17406 162992 76026
rect 163056 19990 163084 79750
rect 163194 79676 163222 80036
rect 163148 79648 163222 79676
rect 163148 79490 163176 79648
rect 163286 79540 163314 80036
rect 163240 79512 163314 79540
rect 163136 79484 163188 79490
rect 163136 79426 163188 79432
rect 163136 78872 163188 78878
rect 163136 78814 163188 78820
rect 163148 77518 163176 78814
rect 163136 77512 163188 77518
rect 163136 77454 163188 77460
rect 163136 76016 163188 76022
rect 163136 75958 163188 75964
rect 163148 21418 163176 75958
rect 163240 21486 163268 79512
rect 163378 79472 163406 80036
rect 163470 79966 163498 80036
rect 163458 79960 163510 79966
rect 163458 79902 163510 79908
rect 163562 79744 163590 80036
rect 163654 79966 163682 80036
rect 163642 79960 163694 79966
rect 163746 79937 163774 80036
rect 163642 79902 163694 79908
rect 163732 79928 163788 79937
rect 163732 79863 163788 79872
rect 163838 79830 163866 80036
rect 163930 79966 163958 80036
rect 164022 79966 164050 80036
rect 164114 79971 164142 80036
rect 163918 79960 163970 79966
rect 163918 79902 163970 79908
rect 164010 79960 164062 79966
rect 164010 79902 164062 79908
rect 164100 79962 164156 79971
rect 164100 79897 164156 79906
rect 163826 79824 163878 79830
rect 163516 79716 163590 79744
rect 163686 79792 163742 79801
rect 164206 79778 164234 80036
rect 164298 79966 164326 80036
rect 164286 79960 164338 79966
rect 164286 79902 164338 79908
rect 163826 79766 163878 79772
rect 163686 79727 163742 79736
rect 164160 79750 164234 79778
rect 163516 79665 163544 79716
rect 163502 79656 163558 79665
rect 163502 79591 163558 79600
rect 163504 79552 163556 79558
rect 163504 79494 163556 79500
rect 163332 79444 163406 79472
rect 163332 49026 163360 79444
rect 163410 78704 163466 78713
rect 163410 78639 163466 78648
rect 163424 76158 163452 78639
rect 163412 76152 163464 76158
rect 163412 76094 163464 76100
rect 163412 75948 163464 75954
rect 163412 75890 163464 75896
rect 163424 71330 163452 75890
rect 163412 71324 163464 71330
rect 163412 71266 163464 71272
rect 163516 70394 163544 79494
rect 163700 75954 163728 79727
rect 163964 79688 164016 79694
rect 164056 79688 164108 79694
rect 163964 79630 164016 79636
rect 164054 79656 164056 79665
rect 164108 79656 164110 79665
rect 163872 79620 163924 79626
rect 163872 79562 163924 79568
rect 163780 79484 163832 79490
rect 163780 79426 163832 79432
rect 163688 75948 163740 75954
rect 163688 75890 163740 75896
rect 163792 75528 163820 79426
rect 163884 76022 163912 79562
rect 163976 76090 164004 79630
rect 164054 79591 164110 79600
rect 164056 78940 164108 78946
rect 164056 78882 164108 78888
rect 164068 77790 164096 78882
rect 164056 77784 164108 77790
rect 164056 77726 164108 77732
rect 163964 76084 164016 76090
rect 163964 76026 164016 76032
rect 163872 76016 163924 76022
rect 163872 75958 163924 75964
rect 163792 75500 163912 75528
rect 163780 75404 163832 75410
rect 163780 75346 163832 75352
rect 163424 70366 163544 70394
rect 163424 64258 163452 70366
rect 163412 64252 163464 64258
rect 163412 64194 163464 64200
rect 163320 49020 163372 49026
rect 163320 48962 163372 48968
rect 163228 21480 163280 21486
rect 163228 21422 163280 21428
rect 163136 21412 163188 21418
rect 163136 21354 163188 21360
rect 163044 19984 163096 19990
rect 163044 19926 163096 19932
rect 162952 17400 163004 17406
rect 162952 17342 163004 17348
rect 162860 13116 162912 13122
rect 162860 13058 162912 13064
rect 162400 11620 162452 11626
rect 162400 11562 162452 11568
rect 161572 10396 161624 10402
rect 161572 10338 161624 10344
rect 161480 6248 161532 6254
rect 161480 6190 161532 6196
rect 162492 4820 162544 4826
rect 162492 4762 162544 4768
rect 161112 4140 161164 4146
rect 161112 4082 161164 4088
rect 161296 3664 161348 3670
rect 161296 3606 161348 3612
rect 161308 480 161336 3606
rect 162504 480 162532 4762
rect 163688 4072 163740 4078
rect 163688 4014 163740 4020
rect 163700 480 163728 4014
rect 163792 3670 163820 75346
rect 163884 75274 163912 75500
rect 164160 75313 164188 79750
rect 164240 79688 164292 79694
rect 164390 79642 164418 80036
rect 164482 79898 164510 80036
rect 164574 79971 164602 80036
rect 164560 79962 164616 79971
rect 164666 79966 164694 80036
rect 164758 79971 164786 80036
rect 164470 79892 164522 79898
rect 164560 79897 164616 79906
rect 164654 79960 164706 79966
rect 164654 79902 164706 79908
rect 164744 79962 164800 79971
rect 164850 79966 164878 80036
rect 164942 79966 164970 80036
rect 165034 79971 165062 80036
rect 164744 79897 164800 79906
rect 164838 79960 164890 79966
rect 164838 79902 164890 79908
rect 164930 79960 164982 79966
rect 164930 79902 164982 79908
rect 165020 79962 165076 79971
rect 165020 79897 165076 79906
rect 164470 79834 164522 79840
rect 164976 79824 165028 79830
rect 164896 79784 164976 79812
rect 164240 79630 164292 79636
rect 164252 78742 164280 79630
rect 164344 79614 164418 79642
rect 164790 79656 164846 79665
rect 164608 79620 164660 79626
rect 164240 78736 164292 78742
rect 164240 78678 164292 78684
rect 164240 77920 164292 77926
rect 164240 77862 164292 77868
rect 164252 76770 164280 77862
rect 164240 76764 164292 76770
rect 164240 76706 164292 76712
rect 164146 75304 164202 75313
rect 163872 75268 163924 75274
rect 164146 75239 164202 75248
rect 163872 75210 163924 75216
rect 164344 11966 164372 79614
rect 164790 79591 164846 79600
rect 164608 79562 164660 79568
rect 164516 79484 164568 79490
rect 164516 79426 164568 79432
rect 164424 78668 164476 78674
rect 164424 78610 164476 78616
rect 164332 11960 164384 11966
rect 164332 11902 164384 11908
rect 164436 11898 164464 78610
rect 164424 11892 164476 11898
rect 164424 11834 164476 11840
rect 164528 11830 164556 79426
rect 164620 78674 164648 79562
rect 164700 79552 164752 79558
rect 164700 79494 164752 79500
rect 164608 78668 164660 78674
rect 164608 78610 164660 78616
rect 164608 78532 164660 78538
rect 164608 78474 164660 78480
rect 164620 76906 164648 78474
rect 164608 76900 164660 76906
rect 164608 76842 164660 76848
rect 164608 75948 164660 75954
rect 164608 75890 164660 75896
rect 164516 11824 164568 11830
rect 164516 11766 164568 11772
rect 164620 11762 164648 75890
rect 164712 14550 164740 79494
rect 164804 17338 164832 79591
rect 164896 75342 164924 79784
rect 165126 79778 165154 80036
rect 165218 79830 165246 80036
rect 165310 79898 165338 80036
rect 165298 79892 165350 79898
rect 165298 79834 165350 79840
rect 164976 79766 165028 79772
rect 165080 79762 165154 79778
rect 165206 79824 165258 79830
rect 165206 79766 165258 79772
rect 165068 79756 165154 79762
rect 165120 79750 165154 79756
rect 165402 79744 165430 80036
rect 165494 79937 165522 80036
rect 165586 79966 165614 80036
rect 165678 79966 165706 80036
rect 165574 79960 165626 79966
rect 165480 79928 165536 79937
rect 165574 79902 165626 79908
rect 165666 79960 165718 79966
rect 165666 79902 165718 79908
rect 165480 79863 165536 79872
rect 165770 79830 165798 80036
rect 165758 79824 165810 79830
rect 165758 79766 165810 79772
rect 165862 79778 165890 80036
rect 165954 79966 165982 80036
rect 165942 79960 165994 79966
rect 166046 79937 166074 80036
rect 165942 79902 165994 79908
rect 166032 79928 166088 79937
rect 166032 79863 166088 79872
rect 165988 79824 166040 79830
rect 165862 79762 165936 79778
rect 165988 79766 166040 79772
rect 166138 79778 166166 80036
rect 166230 79937 166258 80036
rect 166322 79966 166350 80036
rect 166310 79960 166362 79966
rect 166216 79928 166272 79937
rect 166310 79902 166362 79908
rect 166216 79863 166272 79872
rect 166414 79812 166442 80036
rect 166368 79784 166442 79812
rect 165862 79756 165948 79762
rect 165862 79750 165896 79756
rect 165402 79716 165568 79744
rect 165068 79698 165120 79704
rect 164976 79688 165028 79694
rect 164976 79630 165028 79636
rect 165066 79656 165122 79665
rect 164884 75336 164936 75342
rect 164884 75278 164936 75284
rect 164988 71262 165016 79630
rect 165066 79591 165122 79600
rect 165344 79620 165396 79626
rect 164976 71256 165028 71262
rect 164976 71198 165028 71204
rect 165080 70394 165108 79591
rect 165344 79562 165396 79568
rect 165252 79552 165304 79558
rect 165252 79494 165304 79500
rect 165160 79484 165212 79490
rect 165160 79426 165212 79432
rect 165172 76673 165200 79426
rect 165158 76664 165214 76673
rect 165158 76599 165214 76608
rect 165264 75954 165292 79494
rect 165356 75993 165384 79562
rect 165436 79484 165488 79490
rect 165436 79426 165488 79432
rect 165342 75984 165398 75993
rect 165252 75948 165304 75954
rect 165448 75954 165476 79426
rect 165540 78849 165568 79716
rect 165896 79698 165948 79704
rect 165620 79620 165672 79626
rect 165620 79562 165672 79568
rect 165896 79620 165948 79626
rect 165896 79562 165948 79568
rect 165526 78840 165582 78849
rect 165526 78775 165582 78784
rect 165632 78690 165660 79562
rect 165804 79552 165856 79558
rect 165804 79494 165856 79500
rect 165712 78872 165764 78878
rect 165712 78814 165764 78820
rect 165540 78662 165660 78690
rect 165342 75919 165398 75928
rect 165436 75948 165488 75954
rect 165252 75890 165304 75896
rect 165436 75890 165488 75896
rect 165080 70366 165476 70394
rect 164792 17332 164844 17338
rect 164792 17274 164844 17280
rect 164700 14544 164752 14550
rect 164700 14486 164752 14492
rect 164608 11756 164660 11762
rect 164608 11698 164660 11704
rect 165448 9042 165476 70366
rect 165540 17270 165568 78662
rect 165618 77344 165674 77353
rect 165618 77279 165674 77288
rect 165632 76566 165660 77279
rect 165620 76560 165672 76566
rect 165620 76502 165672 76508
rect 165528 17264 165580 17270
rect 165528 17206 165580 17212
rect 165436 9036 165488 9042
rect 165436 8978 165488 8984
rect 165724 8974 165752 78814
rect 165816 76226 165844 79494
rect 165908 77858 165936 79562
rect 166000 79540 166028 79766
rect 166138 79750 166258 79778
rect 166230 79608 166258 79750
rect 166184 79580 166258 79608
rect 166000 79512 166120 79540
rect 165896 77852 165948 77858
rect 165896 77794 165948 77800
rect 165804 76220 165856 76226
rect 165804 76162 165856 76168
rect 165986 75984 166042 75993
rect 165804 75948 165856 75954
rect 165804 75890 165856 75896
rect 165896 75948 165948 75954
rect 165986 75919 166042 75928
rect 165896 75890 165948 75896
rect 165816 14482 165844 75890
rect 165908 22846 165936 75890
rect 166000 22914 166028 75919
rect 166092 22982 166120 79512
rect 166184 78878 166212 79580
rect 166172 78872 166224 78878
rect 166172 78814 166224 78820
rect 166368 78538 166396 79784
rect 166506 79744 166534 80036
rect 166598 79966 166626 80036
rect 166690 79966 166718 80036
rect 166782 79966 166810 80036
rect 166874 79966 166902 80036
rect 166586 79960 166638 79966
rect 166586 79902 166638 79908
rect 166678 79960 166730 79966
rect 166678 79902 166730 79908
rect 166770 79960 166822 79966
rect 166770 79902 166822 79908
rect 166862 79960 166914 79966
rect 166966 79937 166994 80036
rect 166862 79902 166914 79908
rect 166952 79928 167008 79937
rect 166952 79863 167008 79872
rect 167058 79812 167086 80036
rect 167012 79784 167086 79812
rect 166460 79716 166534 79744
rect 166632 79756 166684 79762
rect 166172 78532 166224 78538
rect 166172 78474 166224 78480
rect 166356 78532 166408 78538
rect 166356 78474 166408 78480
rect 166184 31142 166212 78474
rect 166460 78146 166488 79716
rect 166632 79698 166684 79704
rect 166908 79756 166960 79762
rect 166908 79698 166960 79704
rect 166540 79620 166592 79626
rect 166540 79562 166592 79568
rect 166368 78118 166488 78146
rect 166368 75970 166396 78118
rect 166552 76208 166580 79562
rect 166276 75942 166396 75970
rect 166460 76180 166580 76208
rect 166276 65618 166304 75942
rect 166460 71774 166488 76180
rect 166538 75984 166594 75993
rect 166644 75954 166672 79698
rect 166920 79665 166948 79698
rect 166906 79656 166962 79665
rect 166906 79591 166962 79600
rect 167012 79558 167040 79784
rect 167150 79744 167178 80036
rect 167242 79898 167270 80036
rect 167334 79971 167362 80036
rect 167320 79962 167376 79971
rect 167426 79966 167454 80036
rect 167518 79966 167546 80036
rect 167610 79966 167638 80036
rect 167702 79966 167730 80036
rect 167794 79966 167822 80036
rect 167230 79892 167282 79898
rect 167320 79897 167376 79906
rect 167414 79960 167466 79966
rect 167414 79902 167466 79908
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167598 79960 167650 79966
rect 167598 79902 167650 79908
rect 167690 79960 167742 79966
rect 167690 79902 167742 79908
rect 167782 79960 167834 79966
rect 167782 79902 167834 79908
rect 167886 79898 167914 80036
rect 167978 79966 168006 80036
rect 167966 79960 168018 79966
rect 167966 79902 168018 79908
rect 167230 79834 167282 79840
rect 167874 79892 167926 79898
rect 167874 79834 167926 79840
rect 168070 79812 168098 80036
rect 168162 79898 168190 80036
rect 168254 79937 168282 80036
rect 168346 79966 168374 80036
rect 168438 79966 168466 80036
rect 168334 79960 168386 79966
rect 168240 79928 168296 79937
rect 168150 79892 168202 79898
rect 168334 79902 168386 79908
rect 168426 79960 168478 79966
rect 168426 79902 168478 79908
rect 168240 79863 168296 79872
rect 168150 79834 168202 79840
rect 168024 79801 168098 79812
rect 168010 79792 168098 79801
rect 167104 79716 167178 79744
rect 167644 79756 167696 79762
rect 166908 79552 166960 79558
rect 166908 79494 166960 79500
rect 167000 79552 167052 79558
rect 167000 79494 167052 79500
rect 166724 79484 166776 79490
rect 166724 79426 166776 79432
rect 166538 75919 166594 75928
rect 166632 75948 166684 75954
rect 166368 71746 166488 71774
rect 166368 69766 166396 71746
rect 166552 71194 166580 75919
rect 166632 75890 166684 75896
rect 166736 73273 166764 79426
rect 166816 76220 166868 76226
rect 166816 76162 166868 76168
rect 166722 73264 166778 73273
rect 166722 73199 166778 73208
rect 166540 71188 166592 71194
rect 166540 71130 166592 71136
rect 166356 69760 166408 69766
rect 166356 69702 166408 69708
rect 166264 65612 166316 65618
rect 166264 65554 166316 65560
rect 166828 64874 166856 76162
rect 166920 76129 166948 79494
rect 167000 79280 167052 79286
rect 167000 79222 167052 79228
rect 167012 78538 167040 79222
rect 167000 78532 167052 78538
rect 167000 78474 167052 78480
rect 166906 76120 166962 76129
rect 166906 76055 166962 76064
rect 166908 75948 166960 75954
rect 166908 75890 166960 75896
rect 166920 71774 166948 75890
rect 166920 71746 167040 71774
rect 166644 64846 166856 64874
rect 166172 31136 166224 31142
rect 166172 31078 166224 31084
rect 166080 22976 166132 22982
rect 166080 22918 166132 22924
rect 165988 22908 166040 22914
rect 165988 22850 166040 22856
rect 165896 22840 165948 22846
rect 165896 22782 165948 22788
rect 165804 14476 165856 14482
rect 165804 14418 165856 14424
rect 165712 8968 165764 8974
rect 165712 8910 165764 8916
rect 166080 5228 166132 5234
rect 166080 5170 166132 5176
rect 164884 4004 164936 4010
rect 164884 3946 164936 3952
rect 163780 3664 163832 3670
rect 163780 3606 163832 3612
rect 164896 480 164924 3946
rect 166092 480 166120 5170
rect 166644 4826 166672 64846
rect 167012 10334 167040 71746
rect 167104 24478 167132 79716
rect 167644 79698 167696 79704
rect 167736 79756 167788 79762
rect 168066 79784 168098 79792
rect 168288 79824 168340 79830
rect 168380 79824 168432 79830
rect 168288 79766 168340 79772
rect 168378 79792 168380 79801
rect 168432 79792 168434 79801
rect 168010 79727 168066 79736
rect 167736 79698 167788 79704
rect 167460 79688 167512 79694
rect 167512 79648 167592 79676
rect 167460 79630 167512 79636
rect 167276 79620 167328 79626
rect 167276 79562 167328 79568
rect 167368 79620 167420 79626
rect 167368 79562 167420 79568
rect 167184 79484 167236 79490
rect 167184 79426 167236 79432
rect 167092 24472 167144 24478
rect 167092 24414 167144 24420
rect 167196 24274 167224 79426
rect 167288 24410 167316 79562
rect 167380 75954 167408 79562
rect 167460 79552 167512 79558
rect 167460 79494 167512 79500
rect 167472 78878 167500 79494
rect 167460 78872 167512 78878
rect 167460 78814 167512 78820
rect 167368 75948 167420 75954
rect 167368 75890 167420 75896
rect 167460 75948 167512 75954
rect 167460 75890 167512 75896
rect 167368 75744 167420 75750
rect 167368 75686 167420 75692
rect 167276 24404 167328 24410
rect 167276 24346 167328 24352
rect 167380 24342 167408 75686
rect 167472 29646 167500 75890
rect 167564 31074 167592 79648
rect 167656 75750 167684 79698
rect 167748 75954 167776 79698
rect 168104 79688 168156 79694
rect 167932 79648 168104 79676
rect 167828 79620 167880 79626
rect 167828 79562 167880 79568
rect 167736 75948 167788 75954
rect 167736 75890 167788 75896
rect 167644 75744 167696 75750
rect 167644 75686 167696 75692
rect 167840 70394 167868 79562
rect 167932 71058 167960 79648
rect 168104 79630 168156 79636
rect 168196 79688 168248 79694
rect 168196 79630 168248 79636
rect 168102 79520 168158 79529
rect 168102 79455 168158 79464
rect 168012 79280 168064 79286
rect 168012 79222 168064 79228
rect 168024 78606 168052 79222
rect 168116 78713 168144 79455
rect 168102 78704 168158 78713
rect 168102 78639 168158 78648
rect 168012 78600 168064 78606
rect 168012 78542 168064 78548
rect 168208 77489 168236 79630
rect 168194 77480 168250 77489
rect 168194 77415 168250 77424
rect 168010 75984 168066 75993
rect 168010 75919 168066 75928
rect 168024 71126 168052 75919
rect 168300 75177 168328 79766
rect 168530 79744 168558 80036
rect 168378 79727 168434 79736
rect 168484 79716 168558 79744
rect 168380 79552 168432 79558
rect 168380 79494 168432 79500
rect 168286 75168 168342 75177
rect 168286 75103 168342 75112
rect 168012 71120 168064 71126
rect 168012 71062 168064 71068
rect 167920 71052 167972 71058
rect 167920 70994 167972 71000
rect 167656 70366 167868 70394
rect 167656 66978 167684 70366
rect 167644 66972 167696 66978
rect 167644 66914 167696 66920
rect 167552 31068 167604 31074
rect 167552 31010 167604 31016
rect 167460 29640 167512 29646
rect 167460 29582 167512 29588
rect 167368 24336 167420 24342
rect 167368 24278 167420 24284
rect 167184 24268 167236 24274
rect 167184 24210 167236 24216
rect 167000 10328 167052 10334
rect 167000 10270 167052 10276
rect 168392 6186 168420 79494
rect 168484 78810 168512 79716
rect 168622 79676 168650 80036
rect 168714 79898 168742 80036
rect 168806 79971 168834 80036
rect 168792 79962 168848 79971
rect 168898 79966 168926 80036
rect 168990 79971 169018 80036
rect 168702 79892 168754 79898
rect 168792 79897 168848 79906
rect 168886 79960 168938 79966
rect 168886 79902 168938 79908
rect 168976 79962 169032 79971
rect 169082 79966 169110 80036
rect 168976 79897 169032 79906
rect 169070 79960 169122 79966
rect 169070 79902 169122 79908
rect 169174 79898 169202 80036
rect 168702 79834 168754 79840
rect 169162 79892 169214 79898
rect 169162 79834 169214 79840
rect 169266 79830 169294 80036
rect 169358 79830 169386 80036
rect 168932 79824 168984 79830
rect 168932 79766 168984 79772
rect 169024 79824 169076 79830
rect 169024 79766 169076 79772
rect 169254 79824 169306 79830
rect 169254 79766 169306 79772
rect 169346 79824 169398 79830
rect 169450 79801 169478 80036
rect 169542 79966 169570 80036
rect 169530 79960 169582 79966
rect 169530 79902 169582 79908
rect 169634 79898 169662 80036
rect 169726 79898 169754 80036
rect 169818 79898 169846 80036
rect 169910 79937 169938 80036
rect 170002 79966 170030 80036
rect 170094 79966 170122 80036
rect 170186 79966 170214 80036
rect 169990 79960 170042 79966
rect 169896 79928 169952 79937
rect 169622 79892 169674 79898
rect 169622 79834 169674 79840
rect 169714 79892 169766 79898
rect 169714 79834 169766 79840
rect 169806 79892 169858 79898
rect 169990 79902 170042 79908
rect 170082 79960 170134 79966
rect 170082 79902 170134 79908
rect 170174 79960 170226 79966
rect 170174 79902 170226 79908
rect 169896 79863 169952 79872
rect 169806 79834 169858 79840
rect 169944 79824 169996 79830
rect 169346 79766 169398 79772
rect 169436 79792 169492 79801
rect 168576 79648 168650 79676
rect 168746 79656 168802 79665
rect 168472 78804 168524 78810
rect 168472 78746 168524 78752
rect 168576 77194 168604 79648
rect 168746 79591 168802 79600
rect 168840 79620 168892 79626
rect 168656 78804 168708 78810
rect 168656 78746 168708 78752
rect 168484 77166 168604 77194
rect 168484 18698 168512 77166
rect 168564 76492 168616 76498
rect 168564 76434 168616 76440
rect 168472 18692 168524 18698
rect 168472 18634 168524 18640
rect 168576 18630 168604 76434
rect 168668 24206 168696 78746
rect 168760 25770 168788 79591
rect 168840 79562 168892 79568
rect 168852 77194 168880 79562
rect 168944 78810 168972 79766
rect 168932 78804 168984 78810
rect 168932 78746 168984 78752
rect 168852 77166 168972 77194
rect 168840 77104 168892 77110
rect 168840 77046 168892 77052
rect 168852 76974 168880 77046
rect 168840 76968 168892 76974
rect 168840 76910 168892 76916
rect 168944 76498 168972 77166
rect 169036 76498 169064 79766
rect 169116 79756 169168 79762
rect 169850 79792 169906 79801
rect 169436 79727 169492 79736
rect 169576 79756 169628 79762
rect 169116 79698 169168 79704
rect 169576 79698 169628 79704
rect 169668 79756 169720 79762
rect 170278 79812 170306 80036
rect 170370 79966 170398 80036
rect 170462 79971 170490 80036
rect 170358 79960 170410 79966
rect 170358 79902 170410 79908
rect 170448 79962 170504 79971
rect 170554 79966 170582 80036
rect 170646 79966 170674 80036
rect 170448 79897 170504 79906
rect 170542 79960 170594 79966
rect 170542 79902 170594 79908
rect 170634 79960 170686 79966
rect 170634 79902 170686 79908
rect 169944 79766 169996 79772
rect 170232 79784 170306 79812
rect 170496 79824 170548 79830
rect 169850 79727 169906 79736
rect 169668 79698 169720 79704
rect 168932 76492 168984 76498
rect 168932 76434 168984 76440
rect 169024 76492 169076 76498
rect 169024 76434 169076 76440
rect 168840 75132 168892 75138
rect 168840 75074 168892 75080
rect 168748 25764 168800 25770
rect 168748 25706 168800 25712
rect 168852 25702 168880 75074
rect 169128 70394 169156 79698
rect 169390 79656 169446 79665
rect 169208 79620 169260 79626
rect 169208 79562 169260 79568
rect 169312 79614 169390 79642
rect 169220 75138 169248 79562
rect 169208 75132 169260 75138
rect 169208 75074 169260 75080
rect 169312 75002 169340 79614
rect 169390 79591 169446 79600
rect 169484 79620 169536 79626
rect 169484 79562 169536 79568
rect 169392 77988 169444 77994
rect 169392 77930 169444 77936
rect 169404 77450 169432 77930
rect 169392 77444 169444 77450
rect 169392 77386 169444 77392
rect 169300 74996 169352 75002
rect 169300 74938 169352 74944
rect 168944 70366 169156 70394
rect 168944 26926 168972 70366
rect 169496 69698 169524 79562
rect 169588 79370 169616 79698
rect 169680 79665 169708 79698
rect 169760 79688 169812 79694
rect 169666 79656 169722 79665
rect 169760 79630 169812 79636
rect 169666 79591 169722 79600
rect 169588 79342 169708 79370
rect 169576 78736 169628 78742
rect 169576 78678 169628 78684
rect 169588 78130 169616 78678
rect 169576 78124 169628 78130
rect 169576 78066 169628 78072
rect 169680 76537 169708 79342
rect 169666 76528 169722 76537
rect 169666 76463 169722 76472
rect 169772 75206 169800 79630
rect 169864 79558 169892 79727
rect 169852 79552 169904 79558
rect 169852 79494 169904 79500
rect 169956 77976 169984 79766
rect 170036 79688 170088 79694
rect 170036 79630 170088 79636
rect 169864 77948 169984 77976
rect 169760 75200 169812 75206
rect 169760 75142 169812 75148
rect 169760 75064 169812 75070
rect 169760 75006 169812 75012
rect 169484 69692 169536 69698
rect 169484 69634 169536 69640
rect 168932 26920 168984 26926
rect 168932 26862 168984 26868
rect 168840 25696 168892 25702
rect 168840 25638 168892 25644
rect 168656 24200 168708 24206
rect 168656 24142 168708 24148
rect 168564 18624 168616 18630
rect 168564 18566 168616 18572
rect 169772 11665 169800 75006
rect 169864 25634 169892 77948
rect 169942 77480 169998 77489
rect 169942 77415 169998 77424
rect 169956 75546 169984 77415
rect 169944 75540 169996 75546
rect 169944 75482 169996 75488
rect 170048 75426 170076 79630
rect 170128 79620 170180 79626
rect 170128 79562 170180 79568
rect 169956 75398 170076 75426
rect 169852 25628 169904 25634
rect 169852 25570 169904 25576
rect 169956 25566 169984 75398
rect 170036 75200 170088 75206
rect 170036 75142 170088 75148
rect 170048 64190 170076 75142
rect 170140 65550 170168 79562
rect 170232 75070 170260 79784
rect 170496 79766 170548 79772
rect 170404 79756 170456 79762
rect 170404 79698 170456 79704
rect 170312 79552 170364 79558
rect 170312 79494 170364 79500
rect 170324 78742 170352 79494
rect 170312 78736 170364 78742
rect 170312 78678 170364 78684
rect 170416 77353 170444 79698
rect 170508 77489 170536 79766
rect 170588 79756 170640 79762
rect 170588 79698 170640 79704
rect 170600 78062 170628 79698
rect 170738 79676 170766 80036
rect 170830 79801 170858 80036
rect 170816 79792 170872 79801
rect 170816 79727 170872 79736
rect 170922 79676 170950 80036
rect 171014 79744 171042 80036
rect 171106 79937 171134 80036
rect 171198 79966 171226 80036
rect 171186 79960 171238 79966
rect 171092 79928 171148 79937
rect 171186 79902 171238 79908
rect 171092 79863 171148 79872
rect 171290 79812 171318 80036
rect 171382 79971 171410 80036
rect 171368 79962 171424 79971
rect 171368 79897 171424 79906
rect 171290 79784 171364 79812
rect 171014 79716 171088 79744
rect 170738 79648 170812 79676
rect 170922 79648 170996 79676
rect 170588 78056 170640 78062
rect 170588 77998 170640 78004
rect 170784 77994 170812 79648
rect 170772 77988 170824 77994
rect 170772 77930 170824 77936
rect 170588 77852 170640 77858
rect 170588 77794 170640 77800
rect 170494 77480 170550 77489
rect 170494 77415 170550 77424
rect 170402 77344 170458 77353
rect 170402 77279 170458 77288
rect 170312 75540 170364 75546
rect 170312 75482 170364 75488
rect 170220 75064 170272 75070
rect 170220 75006 170272 75012
rect 170324 70394 170352 75482
rect 170600 70394 170628 77794
rect 170680 76560 170732 76566
rect 170680 76502 170732 76508
rect 170232 70366 170352 70394
rect 170508 70366 170628 70394
rect 170232 66910 170260 70366
rect 170220 66904 170272 66910
rect 170220 66846 170272 66852
rect 170128 65544 170180 65550
rect 170128 65486 170180 65492
rect 170036 64184 170088 64190
rect 170036 64126 170088 64132
rect 170508 62830 170536 70366
rect 170496 62824 170548 62830
rect 170496 62766 170548 62772
rect 169944 25560 169996 25566
rect 169944 25502 169996 25508
rect 169758 11656 169814 11665
rect 169758 11591 169814 11600
rect 168380 6180 168432 6186
rect 168380 6122 168432 6128
rect 167184 4956 167236 4962
rect 167184 4898 167236 4904
rect 166632 4820 166684 4826
rect 166632 4762 166684 4768
rect 167196 480 167224 4898
rect 170692 4894 170720 76502
rect 170968 76430 170996 79648
rect 170956 76424 171008 76430
rect 170956 76366 171008 76372
rect 171060 73166 171088 79716
rect 171138 79656 171194 79665
rect 171138 79591 171194 79600
rect 171152 79354 171180 79591
rect 171336 79490 171364 79784
rect 171474 79778 171502 80036
rect 171566 79937 171594 80036
rect 171552 79928 171608 79937
rect 171552 79863 171608 79872
rect 171428 79750 171502 79778
rect 171658 79778 171686 80036
rect 171750 79898 171778 80036
rect 171738 79892 171790 79898
rect 171738 79834 171790 79840
rect 171658 79750 171732 79778
rect 171324 79484 171376 79490
rect 171324 79426 171376 79432
rect 171140 79348 171192 79354
rect 171140 79290 171192 79296
rect 171324 79212 171376 79218
rect 171324 79154 171376 79160
rect 171138 78296 171194 78305
rect 171138 78231 171194 78240
rect 171152 78033 171180 78231
rect 171138 78024 171194 78033
rect 171138 77959 171194 77968
rect 171336 77858 171364 79154
rect 171428 79064 171456 79750
rect 171600 79688 171652 79694
rect 171600 79630 171652 79636
rect 171508 79620 171560 79626
rect 171508 79562 171560 79568
rect 171520 79268 171548 79562
rect 171612 79558 171640 79630
rect 171600 79552 171652 79558
rect 171600 79494 171652 79500
rect 171520 79240 171640 79268
rect 171428 79036 171548 79064
rect 171520 78985 171548 79036
rect 171506 78976 171562 78985
rect 171416 78940 171468 78946
rect 171612 78962 171640 79240
rect 171704 79082 171732 79750
rect 171842 79744 171870 80036
rect 171934 79812 171962 80036
rect 172026 79966 172054 80036
rect 172014 79960 172066 79966
rect 172014 79902 172066 79908
rect 171934 79784 172008 79812
rect 171796 79716 171870 79744
rect 171796 79490 171824 79716
rect 171980 79676 172008 79784
rect 172118 79744 172146 80036
rect 172210 79971 172238 80036
rect 172196 79962 172252 79971
rect 172196 79897 172252 79906
rect 172302 79744 172330 80036
rect 172394 79937 172422 80036
rect 172380 79928 172436 79937
rect 172380 79863 172436 79872
rect 172486 79812 172514 80036
rect 172118 79716 172192 79744
rect 171888 79648 172008 79676
rect 171784 79484 171836 79490
rect 171784 79426 171836 79432
rect 171782 79112 171838 79121
rect 171692 79076 171744 79082
rect 171782 79047 171838 79056
rect 171692 79018 171744 79024
rect 171612 78934 171732 78962
rect 171506 78911 171562 78920
rect 171416 78882 171468 78888
rect 171324 77852 171376 77858
rect 171324 77794 171376 77800
rect 171428 76362 171456 78882
rect 171600 78396 171652 78402
rect 171600 78338 171652 78344
rect 171612 76566 171640 78338
rect 171704 77761 171732 78934
rect 171796 78305 171824 79047
rect 171888 78402 171916 79648
rect 172060 79620 172112 79626
rect 172060 79562 172112 79568
rect 171968 79348 172020 79354
rect 171968 79290 172020 79296
rect 171876 78396 171928 78402
rect 171876 78338 171928 78344
rect 171782 78296 171838 78305
rect 171782 78231 171838 78240
rect 171980 78146 172008 79290
rect 172072 78946 172100 79562
rect 172060 78940 172112 78946
rect 172060 78882 172112 78888
rect 172164 78538 172192 79716
rect 172256 79716 172330 79744
rect 172440 79784 172514 79812
rect 172256 78985 172284 79716
rect 172440 79150 172468 79784
rect 172578 79744 172606 80036
rect 172532 79716 172606 79744
rect 172532 79626 172560 79716
rect 172670 79676 172698 80036
rect 172624 79648 172698 79676
rect 172762 79676 172790 80036
rect 172854 79744 172882 80036
rect 172946 79898 172974 80036
rect 173038 79937 173066 80036
rect 173130 79966 173158 80036
rect 173222 79966 173250 80036
rect 173314 79971 173342 80036
rect 173118 79960 173170 79966
rect 173024 79928 173080 79937
rect 172934 79892 172986 79898
rect 173118 79902 173170 79908
rect 173210 79960 173262 79966
rect 173210 79902 173262 79908
rect 173300 79962 173356 79971
rect 173300 79897 173356 79906
rect 173406 79898 173434 80036
rect 173498 79966 173526 80036
rect 173590 79966 173618 80036
rect 173486 79960 173538 79966
rect 173486 79902 173538 79908
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173024 79863 173080 79872
rect 173394 79892 173446 79898
rect 172934 79834 172986 79840
rect 173394 79834 173446 79840
rect 173072 79824 173124 79830
rect 172978 79792 173034 79801
rect 173072 79766 173124 79772
rect 172854 79716 172928 79744
rect 172978 79727 172980 79736
rect 172762 79648 172836 79676
rect 172520 79620 172572 79626
rect 172520 79562 172572 79568
rect 172518 79520 172574 79529
rect 172518 79455 172574 79464
rect 172532 79354 172560 79455
rect 172520 79348 172572 79354
rect 172520 79290 172572 79296
rect 172336 79144 172388 79150
rect 172336 79086 172388 79092
rect 172428 79144 172480 79150
rect 172428 79086 172480 79092
rect 172242 78976 172298 78985
rect 172242 78911 172298 78920
rect 172152 78532 172204 78538
rect 172152 78474 172204 78480
rect 172060 78464 172112 78470
rect 172060 78406 172112 78412
rect 172072 78282 172100 78406
rect 172072 78254 172192 78282
rect 171980 78118 172100 78146
rect 172072 77926 172100 78118
rect 171968 77920 172020 77926
rect 171968 77862 172020 77868
rect 172060 77920 172112 77926
rect 172060 77862 172112 77868
rect 171690 77752 171746 77761
rect 171690 77687 171746 77696
rect 171784 77716 171836 77722
rect 171784 77658 171836 77664
rect 171692 77648 171744 77654
rect 171692 77590 171744 77596
rect 171600 76560 171652 76566
rect 171600 76502 171652 76508
rect 171416 76356 171468 76362
rect 171416 76298 171468 76304
rect 171048 73160 171100 73166
rect 171048 73102 171100 73108
rect 171140 71528 171192 71534
rect 171140 71470 171192 71476
rect 171152 16574 171180 71470
rect 171704 50386 171732 77590
rect 171796 77364 171824 77658
rect 171796 77336 171916 77364
rect 171784 77104 171836 77110
rect 171784 77046 171836 77052
rect 171796 76770 171824 77046
rect 171784 76764 171836 76770
rect 171784 76706 171836 76712
rect 171888 76650 171916 77336
rect 171796 76622 171916 76650
rect 171692 50380 171744 50386
rect 171692 50322 171744 50328
rect 171796 49094 171824 76622
rect 171876 76560 171928 76566
rect 171876 76502 171928 76508
rect 171784 49088 171836 49094
rect 171784 49030 171836 49036
rect 171152 16546 171824 16574
rect 169576 4888 169628 4894
rect 169576 4830 169628 4836
rect 170680 4888 170732 4894
rect 170680 4830 170732 4836
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 168392 480 168420 3402
rect 169588 480 169616 4830
rect 170772 3528 170824 3534
rect 170772 3470 170824 3476
rect 171796 3482 171824 16546
rect 171888 4078 171916 76502
rect 171980 18834 172008 77862
rect 172060 77580 172112 77586
rect 172060 77522 172112 77528
rect 172072 21622 172100 77522
rect 172164 23118 172192 78254
rect 172244 77784 172296 77790
rect 172244 77726 172296 77732
rect 172256 27062 172284 77726
rect 172348 76770 172376 79086
rect 172428 77852 172480 77858
rect 172428 77794 172480 77800
rect 172336 76764 172388 76770
rect 172336 76706 172388 76712
rect 172336 76356 172388 76362
rect 172336 76298 172388 76304
rect 172244 27056 172296 27062
rect 172244 26998 172296 27004
rect 172152 23112 172204 23118
rect 172152 23054 172204 23060
rect 172060 21616 172112 21622
rect 172060 21558 172112 21564
rect 171968 18828 172020 18834
rect 171968 18770 172020 18776
rect 171876 4072 171928 4078
rect 171876 4014 171928 4020
rect 170784 480 170812 3470
rect 171796 3454 172008 3482
rect 172348 3466 172376 76298
rect 172440 17610 172468 77794
rect 172624 77294 172652 79648
rect 172704 79552 172756 79558
rect 172704 79494 172756 79500
rect 172716 78849 172744 79494
rect 172702 78840 172758 78849
rect 172702 78775 172758 78784
rect 172532 77266 172652 77294
rect 172532 75818 172560 77266
rect 172808 75914 172836 79648
rect 172900 77246 172928 79716
rect 173032 79727 173034 79736
rect 172980 79698 173032 79704
rect 173084 79558 173112 79766
rect 173348 79756 173400 79762
rect 173348 79698 173400 79704
rect 173532 79756 173584 79762
rect 173682 79744 173710 80036
rect 173774 79966 173802 80036
rect 173866 79966 173894 80036
rect 173762 79960 173814 79966
rect 173762 79902 173814 79908
rect 173854 79960 173906 79966
rect 173958 79937 173986 80036
rect 174050 79966 174078 80036
rect 174038 79960 174090 79966
rect 173854 79902 173906 79908
rect 173944 79928 174000 79937
rect 174038 79902 174090 79908
rect 173944 79863 174000 79872
rect 173900 79824 173952 79830
rect 173952 79801 174032 79812
rect 173952 79792 174046 79801
rect 173952 79784 173990 79792
rect 173900 79766 173952 79772
rect 173532 79698 173584 79704
rect 173636 79716 173710 79744
rect 173990 79727 174046 79736
rect 174142 79744 174170 80036
rect 174234 79948 174262 80036
rect 174340 80022 174492 80050
rect 174544 80038 174596 80044
rect 174360 79960 174412 79966
rect 174234 79920 174308 79948
rect 174142 79716 174216 79744
rect 173164 79688 173216 79694
rect 173164 79630 173216 79636
rect 173072 79552 173124 79558
rect 173072 79494 173124 79500
rect 173176 78305 173204 79630
rect 173256 78940 173308 78946
rect 173256 78882 173308 78888
rect 173268 78470 173296 78882
rect 173256 78464 173308 78470
rect 173256 78406 173308 78412
rect 173162 78296 173218 78305
rect 173162 78231 173218 78240
rect 173360 77518 173388 79698
rect 173544 79393 173572 79698
rect 173530 79384 173586 79393
rect 173530 79319 173586 79328
rect 173636 77926 173664 79716
rect 173900 79688 173952 79694
rect 173900 79630 173952 79636
rect 173992 79688 174044 79694
rect 173992 79630 174044 79636
rect 173716 79552 173768 79558
rect 173716 79494 173768 79500
rect 173728 78985 173756 79494
rect 173912 79286 173940 79630
rect 173900 79280 173952 79286
rect 173900 79222 173952 79228
rect 174004 79218 174032 79630
rect 173992 79212 174044 79218
rect 173992 79154 174044 79160
rect 173714 78976 173770 78985
rect 173714 78911 173770 78920
rect 174188 78606 174216 79716
rect 174176 78600 174228 78606
rect 174176 78542 174228 78548
rect 173624 77920 173676 77926
rect 173624 77862 173676 77868
rect 173992 77920 174044 77926
rect 173992 77862 174044 77868
rect 173348 77512 173400 77518
rect 173348 77454 173400 77460
rect 172888 77240 172940 77246
rect 172888 77182 172940 77188
rect 173348 76424 173400 76430
rect 173162 76392 173218 76401
rect 173348 76366 173400 76372
rect 173162 76327 173218 76336
rect 172716 75886 172836 75914
rect 172704 75880 172756 75886
rect 172704 75822 172756 75828
rect 172520 75812 172572 75818
rect 172520 75754 172572 75760
rect 172518 61432 172574 61441
rect 172518 61367 172574 61376
rect 172428 17604 172480 17610
rect 172428 17546 172480 17552
rect 172532 16574 172560 61367
rect 172532 16546 172744 16574
rect 171980 480 172008 3454
rect 172336 3460 172388 3466
rect 172336 3402 172388 3408
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 4010 173204 76327
rect 173254 69592 173310 69601
rect 173254 69527 173310 69536
rect 173164 4004 173216 4010
rect 173164 3946 173216 3952
rect 173268 3534 173296 69527
rect 173360 33114 173388 76366
rect 173898 75712 173954 75721
rect 173898 75647 173954 75656
rect 173348 33108 173400 33114
rect 173348 33050 173400 33056
rect 173256 3528 173308 3534
rect 173256 3470 173308 3476
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 75647
rect 174004 23186 174032 77862
rect 174280 70394 174308 79920
rect 174360 79902 174412 79908
rect 174372 79665 174400 79902
rect 174358 79656 174414 79665
rect 174358 79591 174414 79600
rect 174464 77926 174492 80022
rect 174452 77920 174504 77926
rect 174452 77862 174504 77868
rect 174556 77761 174584 80038
rect 175292 80034 175320 80378
rect 177028 80368 177080 80374
rect 177028 80310 177080 80316
rect 175280 80028 175332 80034
rect 175280 79970 175332 79976
rect 176292 79620 176344 79626
rect 176292 79562 176344 79568
rect 176304 79393 176332 79562
rect 177040 79490 177068 80310
rect 178604 80238 178632 80650
rect 178592 80232 178644 80238
rect 178592 80174 178644 80180
rect 177028 79484 177080 79490
rect 177028 79426 177080 79432
rect 176290 79384 176346 79393
rect 176290 79319 176346 79328
rect 175924 79144 175976 79150
rect 175924 79086 175976 79092
rect 176106 79112 176162 79121
rect 175936 78849 175964 79086
rect 176106 79047 176162 79056
rect 176120 78946 176148 79047
rect 176108 78940 176160 78946
rect 176108 78882 176160 78888
rect 175922 78840 175978 78849
rect 175922 78775 175978 78784
rect 175646 78704 175702 78713
rect 180076 78690 180104 228346
rect 180156 227044 180208 227050
rect 180156 226986 180208 226992
rect 180168 80306 180196 226986
rect 207032 199442 207060 230588
rect 235264 228540 235316 228546
rect 235264 228482 235316 228488
rect 233884 227792 233936 227798
rect 233884 227734 233936 227740
rect 211804 218068 211856 218074
rect 211804 218010 211856 218016
rect 207020 199436 207072 199442
rect 207020 199378 207072 199384
rect 180248 191888 180300 191894
rect 180248 191830 180300 191836
rect 180156 80300 180208 80306
rect 180156 80242 180208 80248
rect 180260 79422 180288 191830
rect 180800 148368 180852 148374
rect 180800 148310 180852 148316
rect 180432 140344 180484 140350
rect 180432 140286 180484 140292
rect 180340 125656 180392 125662
rect 180340 125598 180392 125604
rect 180352 81258 180380 125598
rect 180444 120834 180472 140286
rect 180812 125633 180840 148310
rect 182180 146940 182232 146946
rect 182180 146882 182232 146888
rect 180984 139868 181036 139874
rect 180984 139810 181036 139816
rect 180890 129704 180946 129713
rect 180890 129639 180946 129648
rect 180798 125624 180854 125633
rect 180798 125559 180854 125568
rect 180432 120828 180484 120834
rect 180432 120770 180484 120776
rect 180432 111852 180484 111858
rect 180432 111794 180484 111800
rect 180340 81252 180392 81258
rect 180340 81194 180392 81200
rect 180444 79529 180472 111794
rect 180430 79520 180486 79529
rect 180430 79455 180486 79464
rect 180248 79416 180300 79422
rect 180248 79358 180300 79364
rect 175646 78639 175702 78648
rect 179984 78662 180104 78690
rect 175660 78606 175688 78639
rect 175648 78600 175700 78606
rect 175648 78542 175700 78548
rect 179984 78402 180012 78662
rect 180064 78532 180116 78538
rect 180064 78474 180116 78480
rect 179972 78396 180024 78402
rect 179972 78338 180024 78344
rect 178040 78328 178092 78334
rect 178040 78270 178092 78276
rect 174542 77752 174598 77761
rect 174542 77687 174598 77696
rect 175924 77444 175976 77450
rect 175924 77386 175976 77392
rect 174188 70366 174308 70394
rect 174188 64874 174216 70366
rect 174096 64846 174216 64874
rect 174096 45558 174124 64846
rect 174084 45552 174136 45558
rect 174084 45494 174136 45500
rect 173992 23180 174044 23186
rect 173992 23122 174044 23128
rect 175936 4962 175964 77386
rect 176658 62792 176714 62801
rect 176658 62727 176714 62736
rect 176672 11490 176700 62727
rect 176752 25968 176804 25974
rect 176752 25910 176804 25916
rect 176660 11484 176712 11490
rect 176660 11426 176712 11432
rect 176764 6914 176792 25910
rect 178052 16574 178080 78270
rect 180076 77450 180104 78474
rect 180064 77444 180116 77450
rect 180064 77386 180116 77392
rect 180062 75848 180118 75857
rect 180062 75783 180118 75792
rect 179420 27328 179472 27334
rect 179420 27270 179472 27276
rect 179432 16574 179460 27270
rect 180076 16574 180104 75783
rect 180904 59362 180932 129639
rect 180996 107953 181024 139810
rect 181074 131064 181130 131073
rect 181074 130999 181130 131008
rect 180982 107944 181038 107953
rect 180982 107879 181038 107888
rect 180892 59356 180944 59362
rect 180892 59298 180944 59304
rect 181088 24138 181116 130999
rect 182192 124273 182220 146882
rect 182916 141024 182968 141030
rect 182916 140966 182968 140972
rect 182364 140956 182416 140962
rect 182364 140898 182416 140904
rect 182272 139800 182324 139806
rect 182272 139742 182324 139748
rect 182178 124264 182234 124273
rect 182178 124199 182234 124208
rect 182180 120828 182232 120834
rect 182180 120770 182232 120776
rect 182192 109313 182220 120770
rect 182284 113393 182312 139742
rect 182376 114753 182404 140898
rect 182640 140888 182692 140894
rect 182640 140830 182692 140836
rect 182456 140820 182508 140826
rect 182456 140762 182508 140768
rect 182468 116113 182496 140762
rect 182548 139528 182600 139534
rect 182548 139470 182600 139476
rect 182560 117473 182588 139470
rect 182652 118833 182680 140830
rect 182824 139732 182876 139738
rect 182824 139674 182876 139680
rect 182732 139596 182784 139602
rect 182732 139538 182784 139544
rect 182744 120193 182772 139538
rect 182730 120184 182786 120193
rect 182730 120119 182786 120128
rect 182638 118824 182694 118833
rect 182638 118759 182694 118768
rect 182546 117464 182602 117473
rect 182546 117399 182602 117408
rect 182454 116104 182510 116113
rect 182454 116039 182510 116048
rect 182362 114744 182418 114753
rect 182362 114679 182418 114688
rect 182270 113384 182326 113393
rect 182270 113319 182326 113328
rect 182836 112033 182864 139674
rect 182928 121553 182956 140966
rect 183008 139664 183060 139670
rect 183008 139606 183060 139612
rect 183020 122913 183048 139606
rect 189724 138032 189776 138038
rect 189724 137974 189776 137980
rect 183006 122904 183062 122913
rect 183006 122839 183062 122848
rect 182914 121544 182970 121553
rect 182914 121479 182970 121488
rect 182822 112024 182878 112033
rect 182822 111959 182878 111968
rect 182824 109744 182876 109750
rect 182824 109686 182876 109692
rect 182178 109304 182234 109313
rect 182178 109239 182234 109248
rect 182272 89684 182324 89690
rect 182272 89626 182324 89632
rect 182284 88913 182312 89626
rect 182270 88904 182326 88913
rect 182270 88839 182326 88848
rect 182732 87644 182784 87650
rect 182732 87586 182784 87592
rect 182744 86193 182772 87586
rect 182836 87553 182864 109686
rect 183284 107636 183336 107642
rect 183284 107578 183336 107584
rect 183296 106593 183324 107578
rect 183282 106584 183338 106593
rect 183282 106519 183338 106528
rect 183284 106276 183336 106282
rect 183284 106218 183336 106224
rect 183296 105233 183324 106218
rect 183282 105224 183338 105233
rect 183282 105159 183338 105168
rect 183284 104848 183336 104854
rect 183284 104790 183336 104796
rect 183296 103873 183324 104790
rect 183282 103864 183338 103873
rect 183282 103799 183338 103808
rect 183284 103488 183336 103494
rect 183284 103430 183336 103436
rect 183296 102513 183324 103430
rect 183282 102504 183338 102513
rect 183282 102439 183338 102448
rect 183284 102128 183336 102134
rect 183284 102070 183336 102076
rect 183296 101153 183324 102070
rect 183282 101144 183338 101153
rect 183282 101079 183338 101088
rect 183192 100700 183244 100706
rect 183192 100642 183244 100648
rect 183204 99793 183232 100642
rect 183190 99784 183246 99793
rect 183190 99719 183246 99728
rect 183192 99340 183244 99346
rect 183192 99282 183244 99288
rect 183204 98433 183232 99282
rect 183190 98424 183246 98433
rect 183190 98359 183246 98368
rect 183192 97980 183244 97986
rect 183192 97922 183244 97928
rect 183204 97073 183232 97922
rect 183190 97064 183246 97073
rect 183190 96999 183246 97008
rect 183192 96620 183244 96626
rect 183192 96562 183244 96568
rect 183204 95713 183232 96562
rect 183190 95704 183246 95713
rect 183190 95639 183246 95648
rect 183468 95192 183520 95198
rect 183468 95134 183520 95140
rect 183480 94353 183508 95134
rect 183466 94344 183522 94353
rect 183466 94279 183522 94288
rect 183468 93832 183520 93838
rect 183468 93774 183520 93780
rect 183480 92993 183508 93774
rect 183466 92984 183522 92993
rect 183466 92919 183522 92928
rect 183468 92472 183520 92478
rect 183468 92414 183520 92420
rect 183480 91633 183508 92414
rect 183466 91624 183522 91633
rect 183466 91559 183522 91568
rect 183468 91044 183520 91050
rect 183468 90986 183520 90992
rect 183480 90273 183508 90986
rect 183466 90264 183522 90273
rect 183466 90199 183522 90208
rect 182822 87544 182878 87553
rect 182822 87479 182878 87488
rect 182730 86184 182786 86193
rect 182730 86119 182786 86128
rect 189736 85542 189764 137974
rect 211816 109750 211844 218010
rect 233896 200802 233924 227734
rect 235276 202162 235304 228482
rect 236564 227798 236592 230588
rect 266556 228546 266584 230588
rect 266544 228540 266596 228546
rect 266544 228482 266596 228488
rect 296732 228478 296760 230588
rect 296720 228472 296772 228478
rect 296720 228414 296772 228420
rect 300124 228472 300176 228478
rect 300124 228414 300176 228420
rect 236552 227792 236604 227798
rect 236552 227734 236604 227740
rect 235264 202156 235316 202162
rect 235264 202098 235316 202104
rect 233884 200796 233936 200802
rect 233884 200738 233936 200744
rect 300136 195974 300164 228414
rect 327092 196654 327120 230588
rect 356532 228478 356560 230588
rect 356520 228472 356572 228478
rect 356520 228414 356572 228420
rect 386524 219434 386552 230588
rect 391940 230512 391992 230518
rect 391940 230454 391992 230460
rect 391952 223582 391980 230454
rect 389824 223576 389876 223582
rect 389824 223518 389876 223524
rect 391940 223576 391992 223582
rect 391940 223518 391992 223524
rect 386432 219406 386552 219434
rect 378324 214600 378376 214606
rect 378324 214542 378376 214548
rect 378336 212566 378364 214542
rect 378324 212560 378376 212566
rect 378324 212502 378376 212508
rect 374920 212492 374972 212498
rect 374920 212434 374972 212440
rect 374932 209846 374960 212434
rect 370504 209840 370556 209846
rect 370504 209782 370556 209788
rect 374920 209840 374972 209846
rect 374920 209782 374972 209788
rect 370516 197402 370544 209782
rect 386432 198014 386460 219406
rect 389836 218142 389864 223518
rect 387800 218136 387852 218142
rect 387800 218078 387852 218084
rect 389824 218136 389876 218142
rect 389824 218078 389876 218084
rect 387812 214606 387840 218078
rect 387800 214600 387852 214606
rect 387800 214542 387852 214548
rect 386420 198008 386472 198014
rect 386420 197950 386472 197956
rect 367744 197396 367796 197402
rect 367744 197338 367796 197344
rect 370504 197396 370556 197402
rect 370504 197338 370556 197344
rect 327080 196648 327132 196654
rect 327080 196590 327132 196596
rect 300124 195968 300176 195974
rect 300124 195910 300176 195916
rect 211896 178084 211948 178090
rect 211896 178026 211948 178032
rect 211804 109744 211856 109750
rect 211804 109686 211856 109692
rect 211908 87650 211936 178026
rect 367756 176730 367784 197338
rect 366364 176724 366416 176730
rect 366364 176666 366416 176672
rect 367744 176724 367796 176730
rect 367744 176666 367796 176672
rect 345664 151836 345716 151842
rect 345664 151778 345716 151784
rect 238024 99408 238076 99414
rect 238024 99350 238076 99356
rect 211896 87644 211948 87650
rect 211896 87586 211948 87592
rect 182732 85536 182784 85542
rect 182732 85478 182784 85484
rect 189724 85536 189776 85542
rect 189724 85478 189776 85484
rect 182744 84833 182772 85478
rect 182730 84824 182786 84833
rect 182730 84759 182786 84768
rect 238036 84182 238064 99350
rect 182732 84176 182784 84182
rect 182732 84118 182784 84124
rect 238024 84176 238076 84182
rect 238024 84118 238076 84124
rect 182744 83473 182772 84118
rect 182730 83464 182786 83473
rect 182730 83399 182786 83408
rect 182914 82104 182970 82113
rect 182914 82039 182970 82048
rect 182822 80744 182878 80753
rect 182822 80679 182878 80688
rect 182836 24138 182864 80679
rect 182928 60722 182956 82039
rect 345676 80782 345704 151778
rect 366376 138106 366404 176666
rect 361580 138100 361632 138106
rect 361580 138042 361632 138048
rect 366364 138100 366416 138106
rect 366364 138042 366416 138048
rect 361592 135318 361620 138042
rect 360844 135312 360896 135318
rect 360844 135254 360896 135260
rect 361580 135312 361632 135318
rect 361580 135254 361632 135260
rect 360856 131170 360884 135254
rect 359464 131164 359516 131170
rect 359464 131106 359516 131112
rect 360844 131164 360896 131170
rect 360844 131106 360896 131112
rect 359476 110498 359504 131106
rect 357440 110492 357492 110498
rect 357440 110434 357492 110440
rect 359464 110492 359516 110498
rect 359464 110434 359516 110440
rect 357452 107642 357480 110434
rect 357440 107636 357492 107642
rect 357440 107578 357492 107584
rect 345664 80776 345716 80782
rect 345664 80718 345716 80724
rect 393976 80617 394004 231814
rect 394804 230518 394832 232222
rect 394792 230512 394844 230518
rect 394792 230454 394844 230460
rect 396460 106282 396488 700334
rect 396724 643136 396776 643142
rect 396724 643078 396776 643084
rect 396540 411936 396592 411942
rect 396540 411878 396592 411884
rect 396552 232286 396580 411878
rect 396540 232280 396592 232286
rect 396540 232222 396592 232228
rect 396448 106276 396500 106282
rect 396448 106218 396500 106224
rect 393962 80608 394018 80617
rect 393962 80543 394018 80552
rect 356060 80232 356112 80238
rect 356060 80174 356112 80180
rect 242164 78260 242216 78266
rect 242164 78202 242216 78208
rect 226340 77172 226392 77178
rect 226340 77114 226392 77120
rect 190460 76492 190512 76498
rect 190460 76434 190512 76440
rect 184940 68468 184992 68474
rect 184940 68410 184992 68416
rect 182916 60716 182968 60722
rect 182916 60658 182968 60664
rect 183560 27260 183612 27266
rect 183560 27202 183612 27208
rect 181076 24132 181128 24138
rect 181076 24074 181128 24080
rect 182824 24132 182876 24138
rect 182824 24074 182876 24080
rect 183572 16574 183600 27202
rect 178052 16546 178632 16574
rect 179432 16546 180012 16574
rect 180076 16546 180380 16574
rect 183572 16546 183784 16574
rect 177856 11484 177908 11490
rect 177856 11426 177908 11432
rect 176672 6886 176792 6914
rect 175924 4956 175976 4962
rect 175924 4898 175976 4904
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 175476 480 175504 3470
rect 176672 480 176700 6886
rect 177868 480 177896 11426
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 179984 3482 180012 16546
rect 179984 3454 180288 3482
rect 180352 3466 180380 16546
rect 181444 6860 181496 6866
rect 181444 6802 181496 6808
rect 180260 480 180288 3454
rect 180340 3460 180392 3466
rect 180340 3402 180392 3408
rect 181456 480 181484 6802
rect 182548 4140 182600 4146
rect 182548 4082 182600 4088
rect 182560 480 182588 4082
rect 183756 480 183784 16546
rect 184952 11558 184980 68410
rect 189080 67108 189132 67114
rect 189080 67050 189132 67056
rect 186320 27192 186372 27198
rect 186320 27134 186372 27140
rect 186332 16574 186360 27134
rect 189092 16574 189120 67050
rect 186332 16546 186912 16574
rect 189092 16546 189304 16574
rect 184940 11552 184992 11558
rect 184940 11494 184992 11500
rect 186136 11552 186188 11558
rect 186136 11494 186188 11500
rect 184940 11416 184992 11422
rect 184940 11358 184992 11364
rect 184952 480 184980 11358
rect 186148 480 186176 11494
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188528 14340 188580 14346
rect 188528 14282 188580 14288
rect 188540 480 188568 14282
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 76434
rect 194598 75576 194654 75585
rect 194598 75511 194654 75520
rect 193218 65512 193274 65521
rect 193218 65447 193274 65456
rect 191838 17096 191894 17105
rect 191838 17031 191894 17040
rect 191852 16574 191880 17031
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 65447
rect 194612 16574 194640 75511
rect 209780 73976 209832 73982
rect 209780 73918 209832 73924
rect 198740 32904 198792 32910
rect 198740 32846 198792 32852
rect 194612 16546 195192 16574
rect 194414 6080 194470 6089
rect 194414 6015 194470 6024
rect 194428 480 194456 6015
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 197910 8800 197966 8809
rect 197910 8735 197966 8744
rect 196808 4072 196860 4078
rect 196808 4014 196860 4020
rect 196820 480 196848 4014
rect 197924 480 197952 8735
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 32846
rect 201500 32836 201552 32842
rect 201500 32778 201552 32784
rect 201512 11558 201540 32778
rect 201592 28620 201644 28626
rect 201592 28562 201644 28568
rect 201500 11552 201552 11558
rect 201500 11494 201552 11500
rect 201604 6914 201632 28562
rect 204260 28552 204312 28558
rect 204260 28494 204312 28500
rect 204272 16574 204300 28494
rect 208400 28484 208452 28490
rect 208400 28426 208452 28432
rect 208412 16574 208440 28426
rect 204272 16546 205128 16574
rect 208412 16546 208624 16574
rect 202696 11552 202748 11558
rect 202696 11494 202748 11500
rect 201512 6886 201632 6914
rect 200304 3936 200356 3942
rect 200304 3878 200356 3884
rect 200316 480 200344 3878
rect 201512 480 201540 6886
rect 202708 480 202736 11494
rect 203892 3868 203944 3874
rect 203892 3810 203944 3816
rect 203904 480 203932 3810
rect 205100 480 205128 16546
rect 206192 5160 206244 5166
rect 206192 5102 206244 5108
rect 206204 480 206232 5102
rect 207388 3596 207440 3602
rect 207388 3538 207440 3544
rect 207400 480 207428 3538
rect 208596 480 208624 16546
rect 209792 480 209820 73918
rect 223580 73908 223632 73914
rect 223580 73850 223632 73856
rect 218704 68400 218756 68406
rect 218704 68342 218756 68348
rect 212538 34096 212594 34105
rect 212538 34031 212594 34040
rect 212552 16574 212580 34031
rect 215300 29980 215352 29986
rect 215300 29922 215352 29928
rect 212552 16546 213408 16574
rect 210974 4040 211030 4049
rect 210974 3975 211030 3984
rect 212172 4004 212224 4010
rect 210988 480 211016 3975
rect 212172 3946 212224 3952
rect 212184 480 212212 3946
rect 213380 480 213408 16546
rect 214470 3224 214526 3233
rect 214470 3159 214526 3168
rect 214484 480 214512 3159
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 29922
rect 218060 27124 218112 27130
rect 218060 27066 218112 27072
rect 216680 17876 216732 17882
rect 216680 17818 216732 17824
rect 216692 16574 216720 17818
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 3602 218100 27066
rect 218716 4146 218744 68342
rect 219440 33856 219492 33862
rect 219440 33798 219492 33804
rect 219452 16574 219480 33798
rect 219452 16546 220032 16574
rect 218704 4140 218756 4146
rect 218704 4082 218756 4088
rect 219348 4140 219400 4146
rect 219348 4082 219400 4088
rect 218150 3904 218206 3913
rect 218150 3839 218206 3848
rect 218060 3596 218112 3602
rect 218060 3538 218112 3544
rect 218164 1986 218192 3839
rect 219360 3602 219388 4082
rect 219256 3596 219308 3602
rect 219256 3538 219308 3544
rect 219348 3596 219400 3602
rect 219348 3538 219400 3544
rect 218072 1958 218192 1986
rect 218072 480 218100 1958
rect 219268 480 219296 3538
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 222752 7880 222804 7886
rect 222752 7822 222804 7828
rect 221554 3768 221610 3777
rect 221554 3703 221610 3712
rect 221568 480 221596 3703
rect 222764 480 222792 7822
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 73850
rect 224960 63028 225012 63034
rect 224960 62970 225012 62976
rect 224972 16574 225000 62970
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 77114
rect 230478 74080 230534 74089
rect 230478 74015 230534 74024
rect 226430 33960 226486 33969
rect 226430 33895 226486 33904
rect 226444 16574 226472 33895
rect 230492 16574 230520 74015
rect 234620 33788 234672 33794
rect 234620 33730 234672 33736
rect 226444 16546 227576 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 229374 13288 229430 13297
rect 229374 13223 229430 13232
rect 228730 6896 228786 6905
rect 228730 6831 228786 6840
rect 228744 480 228772 6831
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 13223
rect 231044 480 231072 16546
rect 233424 11688 233476 11694
rect 233424 11630 233476 11636
rect 232228 3800 232280 3806
rect 232228 3742 232280 3748
rect 232240 480 232268 3742
rect 233436 480 233464 11630
rect 234632 480 234660 33730
rect 242176 20466 242204 78202
rect 304264 78192 304316 78198
rect 255962 78160 256018 78169
rect 304264 78134 304316 78140
rect 255962 78095 256018 78104
rect 249800 77104 249852 77110
rect 249800 77046 249852 77052
rect 247040 77036 247092 77042
rect 247040 76978 247092 76984
rect 244278 73944 244334 73953
rect 244278 73879 244334 73888
rect 242898 27024 242954 27033
rect 242898 26959 242954 26968
rect 242164 20460 242216 20466
rect 242164 20402 242216 20408
rect 241520 18896 241572 18902
rect 241520 18838 241572 18844
rect 241532 16574 241560 18838
rect 241532 16546 241744 16574
rect 237656 16244 237708 16250
rect 237656 16186 237708 16192
rect 236552 12436 236604 12442
rect 236552 12378 236604 12384
rect 235814 3632 235870 3641
rect 235814 3567 235870 3576
rect 235828 480 235856 3567
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 12378
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16186
rect 240140 11620 240192 11626
rect 240140 11562 240192 11568
rect 239312 6792 239364 6798
rect 239312 6734 239364 6740
rect 239324 480 239352 6734
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 11562
rect 241716 480 241744 16546
rect 242912 3398 242940 26959
rect 244292 16574 244320 73879
rect 247052 16574 247080 76978
rect 248418 20496 248474 20505
rect 248418 20431 248474 20440
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 242992 6724 243044 6730
rect 242992 6666 243044 6672
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 243004 3210 243032 6666
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242912 3182 243032 3210
rect 242912 480 242940 3182
rect 244108 480 244136 3334
rect 245212 480 245240 16546
rect 246394 6760 246450 6769
rect 246394 6695 246450 6704
rect 246408 480 246436 6695
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 20431
rect 249812 16574 249840 77046
rect 255976 20534 256004 78095
rect 282918 77208 282974 77217
rect 282918 77143 282974 77152
rect 260840 76968 260892 76974
rect 260840 76910 260892 76916
rect 255320 20528 255372 20534
rect 255320 20470 255372 20476
rect 255964 20528 256016 20534
rect 255964 20470 256016 20476
rect 251178 17912 251234 17921
rect 251178 17847 251234 17856
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3806 251220 17847
rect 255332 16574 255360 20470
rect 259460 19916 259512 19922
rect 259460 19858 259512 19864
rect 255332 16546 255912 16574
rect 254216 15156 254268 15162
rect 254216 15098 254268 15104
rect 251272 14408 251324 14414
rect 251272 14350 251324 14356
rect 251180 3800 251232 3806
rect 251180 3742 251232 3748
rect 251284 3482 251312 14350
rect 253480 6656 253532 6662
rect 253480 6598 253532 6604
rect 252376 3800 252428 3806
rect 252376 3742 252428 3748
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3742
rect 253492 480 253520 6598
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 15098
rect 255884 480 255912 16546
rect 258264 15088 258316 15094
rect 258264 15030 258316 15036
rect 257068 6588 257120 6594
rect 257068 6530 257120 6536
rect 257080 480 257108 6530
rect 258276 480 258304 15030
rect 259472 480 259500 19858
rect 260852 16574 260880 76910
rect 266358 33824 266414 33833
rect 266358 33759 266414 33768
rect 262220 20664 262272 20670
rect 262220 20606 262272 20612
rect 262232 16574 262260 20606
rect 266372 16574 266400 33759
rect 269120 17808 269172 17814
rect 269120 17750 269172 17756
rect 280158 17776 280214 17785
rect 269132 16574 269160 17750
rect 273260 17740 273312 17746
rect 280158 17711 280214 17720
rect 273260 17682 273312 17688
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 260656 6520 260708 6526
rect 260656 6462 260708 6468
rect 260668 480 260696 6462
rect 261772 480 261800 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264978 14920 265034 14929
rect 264978 14855 265034 14864
rect 264150 6624 264206 6633
rect 264150 6559 264206 6568
rect 264164 480 264192 6559
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 14855
rect 266556 480 266584 16546
rect 268384 15020 268436 15026
rect 268384 14962 268436 14968
rect 267740 3732 267792 3738
rect 267740 3674 267792 3680
rect 267752 480 267780 3674
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 14962
rect 270052 480 270080 16546
rect 272432 14952 272484 14958
rect 272432 14894 272484 14900
rect 271236 6452 271288 6458
rect 271236 6394 271288 6400
rect 271248 480 271276 6394
rect 272444 480 272472 14894
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 17682
rect 276020 17672 276072 17678
rect 276020 17614 276072 17620
rect 274824 6384 274876 6390
rect 274824 6326 274876 6332
rect 274836 480 274864 6326
rect 276032 3738 276060 17614
rect 280172 16574 280200 17711
rect 282932 16574 282960 77143
rect 284300 76900 284352 76906
rect 284300 76842 284352 76848
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 279054 14784 279110 14793
rect 279054 14719 279110 14728
rect 276112 12368 276164 12374
rect 276112 12310 276164 12316
rect 276020 3732 276072 3738
rect 276020 3674 276072 3680
rect 276124 3482 276152 12310
rect 278320 9580 278372 9586
rect 278320 9522 278372 9528
rect 276756 3732 276808 3738
rect 276756 3674 276808 3680
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3674
rect 278332 480 278360 9522
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 14719
rect 280724 480 280752 16546
rect 281906 9616 281962 9625
rect 281906 9551 281962 9560
rect 281920 480 281948 9551
rect 283116 480 283144 16546
rect 284312 3738 284340 76842
rect 296720 76832 296772 76838
rect 296720 76774 296772 76780
rect 291200 35420 291252 35426
rect 291200 35362 291252 35368
rect 285680 32768 285732 32774
rect 285680 32710 285732 32716
rect 284390 17640 284446 17649
rect 284390 17575 284446 17584
rect 284300 3732 284352 3738
rect 284300 3674 284352 3680
rect 284404 3482 284432 17575
rect 285692 16574 285720 32710
rect 287060 32700 287112 32706
rect 287060 32642 287112 32648
rect 287072 16574 287100 32642
rect 289820 25900 289872 25906
rect 289820 25842 289872 25848
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 285036 3732 285088 3738
rect 285036 3674 285088 3680
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3674
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288992 9512 289044 9518
rect 288992 9454 289044 9460
rect 289004 480 289032 9454
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 25842
rect 291212 16574 291240 35362
rect 292580 24540 292632 24546
rect 292580 24482 292632 24488
rect 292592 16574 292620 24482
rect 296732 16574 296760 76774
rect 298098 72584 298154 72593
rect 298098 72519 298154 72528
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 296732 16546 297312 16574
rect 291396 480 291424 16546
rect 292580 9444 292632 9450
rect 292580 9386 292632 9392
rect 292592 480 292620 9386
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 296076 9376 296128 9382
rect 296076 9318 296128 9324
rect 294880 5092 294932 5098
rect 294880 5034 294932 5040
rect 294892 480 294920 5034
rect 296088 480 296116 9318
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 72519
rect 303620 61464 303672 61470
rect 303620 61406 303672 61412
rect 300858 17504 300914 17513
rect 300858 17439 300914 17448
rect 300872 16574 300900 17439
rect 303632 16574 303660 61406
rect 304276 31210 304304 78134
rect 354678 77072 354734 77081
rect 354678 77007 354734 77016
rect 318800 73840 318852 73846
rect 318800 73782 318852 73788
rect 305000 72820 305052 72826
rect 305000 72762 305052 72768
rect 304264 31204 304316 31210
rect 304264 31146 304316 31152
rect 305012 16574 305040 72762
rect 307760 72752 307812 72758
rect 307760 72694 307812 72700
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299662 9480 299718 9489
rect 299662 9415 299718 9424
rect 299676 480 299704 9415
rect 300766 6488 300822 6497
rect 300766 6423 300822 6432
rect 300780 480 300808 6423
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303160 9308 303212 9314
rect 303160 9250 303212 9256
rect 303172 480 303200 9250
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 9240 306800 9246
rect 306748 9182 306800 9188
rect 306760 480 306788 9182
rect 307772 3398 307800 72694
rect 311900 72684 311952 72690
rect 311900 72626 311952 72632
rect 311912 16574 311940 72626
rect 316038 35320 316094 35329
rect 316038 35255 316094 35264
rect 316052 16574 316080 35255
rect 317418 26888 317474 26897
rect 317418 26823 317474 26832
rect 317432 16574 317460 26823
rect 318812 16574 318840 73782
rect 332600 72616 332652 72622
rect 332600 72558 332652 72564
rect 320180 68332 320232 68338
rect 320180 68274 320232 68280
rect 320192 16574 320220 68274
rect 331220 60240 331272 60246
rect 331220 60182 331272 60188
rect 325700 57316 325752 57322
rect 325700 57258 325752 57264
rect 321560 32632 321612 32638
rect 321560 32574 321612 32580
rect 321572 16574 321600 32574
rect 325712 16574 325740 57258
rect 329840 20596 329892 20602
rect 329840 20538 329892 20544
rect 329852 16574 329880 20538
rect 311912 16546 312216 16574
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 325712 16546 326384 16574
rect 329852 16546 330432 16574
rect 311440 14884 311492 14890
rect 311440 14826 311492 14832
rect 310244 9172 310296 9178
rect 310244 9114 310296 9120
rect 307944 7812 307996 7818
rect 307944 7754 307996 7760
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 7754
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 9114
rect 311452 480 311480 14826
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 315026 9344 315082 9353
rect 315026 9279 315082 9288
rect 313832 9104 313884 9110
rect 313832 9046 313884 9052
rect 313844 480 313872 9046
rect 315040 480 315068 9279
rect 316236 480 316264 16546
rect 317326 9208 317382 9217
rect 317326 9143 317382 9152
rect 317340 480 317368 9143
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 324412 10464 324464 10470
rect 324412 10406 324464 10412
rect 323308 7744 323360 7750
rect 323308 7686 323360 7692
rect 323320 480 323348 7686
rect 324320 3664 324372 3670
rect 324320 3606 324372 3612
rect 324332 1850 324360 3606
rect 324424 3398 324452 10406
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 1822 324452 1850
rect 324424 480 324452 1822
rect 325620 480 325648 3334
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328000 12300 328052 12306
rect 328000 12242 328052 12248
rect 328012 480 328040 12242
rect 328736 12232 328788 12238
rect 328736 12174 328788 12180
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 12174
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 60182
rect 332612 3398 332640 72558
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 338120 64524 338172 64530
rect 338120 64466 338172 64472
rect 336738 31104 336794 31113
rect 336738 31039 336794 31048
rect 332692 28416 332744 28422
rect 332692 28358 332744 28364
rect 335358 28384 335414 28393
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 28358
rect 335358 28319 335414 28328
rect 335372 16574 335400 28319
rect 336752 16574 336780 31039
rect 338132 16574 338160 64466
rect 339500 64456 339552 64462
rect 339500 64398 339552 64404
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 334622 12064 334678 12073
rect 334622 11999 334678 12008
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 11999
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 64398
rect 340892 3210 340920 72490
rect 353298 68232 353354 68241
rect 353298 68167 353354 68176
rect 340972 62960 341024 62966
rect 340972 62902 341024 62908
rect 340984 3398 341012 62902
rect 351918 51776 351974 51785
rect 351918 51711 351974 51720
rect 346400 32564 346452 32570
rect 346400 32506 346452 32512
rect 343640 21684 343692 21690
rect 343640 21626 343692 21632
rect 343652 16574 343680 21626
rect 346412 16574 346440 32506
rect 349160 32496 349212 32502
rect 349160 32438 349212 32444
rect 347780 17604 347832 17610
rect 347780 17546 347832 17552
rect 347792 16574 347820 17546
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 342904 16176 342956 16182
rect 342904 16118 342956 16124
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16118
rect 344572 480 344600 16546
rect 345296 12164 345348 12170
rect 345296 12106 345348 12112
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 12106
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 1562 349200 32438
rect 351932 16574 351960 51711
rect 353312 16574 353340 68167
rect 354692 16574 354720 77007
rect 356072 16574 356100 80174
rect 374000 80164 374052 80170
rect 374000 80106 374052 80112
rect 368480 72480 368532 72486
rect 368480 72422 368532 72428
rect 367100 65680 367152 65686
rect 367100 65622 367152 65628
rect 362960 60172 363012 60178
rect 362960 60114 363012 60120
rect 357440 50448 357492 50454
rect 357440 50390 357492 50396
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349252 13456 349304 13462
rect 349252 13398 349304 13404
rect 349160 1556 349212 1562
rect 349160 1498 349212 1504
rect 349264 480 349292 13398
rect 351642 9072 351698 9081
rect 351642 9007 351698 9016
rect 350448 1556 350500 1562
rect 350448 1498 350500 1504
rect 350460 480 350488 1498
rect 351656 480 351684 9007
rect 352852 480 352880 16546
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3398 357480 50390
rect 362972 16574 363000 60114
rect 367112 16574 367140 65622
rect 368492 16574 368520 72422
rect 372618 58576 372674 58585
rect 372618 58511 372674 58520
rect 372632 16574 372660 58511
rect 362972 16546 363552 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 372632 16546 372936 16574
rect 361120 16108 361172 16114
rect 361120 16050 361172 16056
rect 357532 13388 357584 13394
rect 357532 13330 357584 13336
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 13330
rect 359464 13320 359516 13326
rect 359464 13262 359516 13268
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 13262
rect 361132 480 361160 16050
rect 361856 13252 361908 13258
rect 361856 13194 361908 13200
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 13194
rect 363524 480 363552 16546
rect 365718 16144 365774 16153
rect 365718 16079 365774 16088
rect 364616 5024 364668 5030
rect 364616 4966 364668 4972
rect 364628 480 364656 4966
rect 365732 3210 365760 16079
rect 365812 13184 365864 13190
rect 365812 13126 365864 13132
rect 365824 3398 365852 13126
rect 365812 3392 365864 3398
rect 365812 3334 365864 3340
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 365732 3182 365852 3210
rect 365824 480 365852 3182
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 370134 14648 370190 14657
rect 370134 14583 370190 14592
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 14583
rect 371238 13152 371294 13161
rect 371238 13087 371294 13096
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 13087
rect 372908 480 372936 16546
rect 374012 1170 374040 80106
rect 396736 77450 396764 643078
rect 396816 404388 396868 404394
rect 396816 404330 396868 404336
rect 396828 142866 396856 404330
rect 396908 351960 396960 351966
rect 396908 351902 396960 351908
rect 396816 142860 396868 142866
rect 396816 142802 396868 142808
rect 396920 140214 396948 351902
rect 397000 298172 397052 298178
rect 397000 298114 397052 298120
rect 397012 140282 397040 298114
rect 397092 244316 397144 244322
rect 397092 244258 397144 244264
rect 397104 141778 397132 244258
rect 397092 141772 397144 141778
rect 397092 141714 397144 141720
rect 397000 140276 397052 140282
rect 397000 140218 397052 140224
rect 396908 140208 396960 140214
rect 396908 140150 396960 140156
rect 397472 78849 397500 703520
rect 413664 700466 413692 703520
rect 397644 700460 397696 700466
rect 397644 700402 397696 700408
rect 405004 700460 405056 700466
rect 405004 700402 405056 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 397552 700324 397604 700330
rect 397552 700266 397604 700272
rect 397458 78840 397514 78849
rect 397458 78775 397514 78784
rect 397564 78538 397592 700266
rect 397656 231130 397684 700402
rect 403624 700392 403676 700398
rect 403624 700334 403676 700340
rect 400864 700324 400916 700330
rect 400864 700266 400916 700272
rect 398104 696992 398156 696998
rect 398104 696934 398156 696940
rect 397644 231124 397696 231130
rect 397644 231066 397696 231072
rect 398116 78674 398144 696934
rect 399484 683188 399536 683194
rect 399484 683130 399536 683136
rect 398196 378208 398248 378214
rect 398196 378150 398248 378156
rect 398208 79082 398236 378150
rect 399496 100706 399524 683130
rect 400876 102134 400904 700266
rect 403636 103494 403664 700334
rect 405016 104854 405044 700402
rect 417424 630692 417476 630698
rect 417424 630634 417476 630640
rect 414664 576904 414716 576910
rect 414664 576846 414716 576852
rect 413284 524476 413336 524482
rect 413284 524418 413336 524424
rect 409144 418192 409196 418198
rect 409144 418134 409196 418140
rect 407764 311908 407816 311914
rect 407764 311850 407816 311856
rect 406384 258120 406436 258126
rect 406384 258062 406436 258068
rect 405004 104848 405056 104854
rect 405004 104790 405056 104796
rect 403624 103488 403676 103494
rect 403624 103430 403676 103436
rect 400864 102128 400916 102134
rect 400864 102070 400916 102076
rect 399484 100700 399536 100706
rect 399484 100642 399536 100648
rect 406396 89690 406424 258062
rect 407776 91050 407804 311850
rect 409156 93838 409184 418134
rect 413296 96626 413324 524418
rect 414676 97986 414704 576846
rect 417436 99346 417464 630634
rect 418804 364404 418856 364410
rect 418804 364346 418856 364352
rect 417424 99340 417476 99346
rect 417424 99282 417476 99288
rect 414664 97980 414716 97986
rect 414664 97922 414716 97928
rect 413284 96620 413336 96626
rect 413284 96562 413336 96568
rect 409144 93832 409196 93838
rect 409144 93774 409196 93780
rect 418816 92478 418844 364346
rect 429212 141710 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 141704 429252 141710
rect 429200 141646 429252 141652
rect 418804 92472 418856 92478
rect 418804 92414 418856 92420
rect 407764 91044 407816 91050
rect 407764 90986 407816 90992
rect 406384 89684 406436 89690
rect 406384 89626 406436 89632
rect 426440 80096 426492 80102
rect 426440 80038 426492 80044
rect 398196 79076 398248 79082
rect 398196 79018 398248 79024
rect 398104 78668 398156 78674
rect 398104 78610 398156 78616
rect 397552 78532 397604 78538
rect 397552 78474 397604 78480
rect 396724 77444 396776 77450
rect 396724 77386 396776 77392
rect 389178 76936 389234 76945
rect 389178 76871 389234 76880
rect 376760 76764 376812 76770
rect 376760 76706 376812 76712
rect 375380 76696 375432 76702
rect 375380 76638 375432 76644
rect 374092 58744 374144 58750
rect 374092 58686 374144 58692
rect 374104 3398 374132 58686
rect 375392 16574 375420 76638
rect 376772 16574 376800 76706
rect 382280 71460 382332 71466
rect 382280 71402 382332 71408
rect 378140 28348 378192 28354
rect 378140 28290 378192 28296
rect 378152 16574 378180 28290
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379520 14816 379572 14822
rect 379520 14758 379572 14764
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 14758
rect 381176 14748 381228 14754
rect 381176 14690 381228 14696
rect 381188 480 381216 14690
rect 382292 3210 382320 71402
rect 382372 35352 382424 35358
rect 382372 35294 382424 35300
rect 382384 3398 382412 35294
rect 389192 16574 389220 76871
rect 402978 75440 403034 75449
rect 402978 75375 403034 75384
rect 390560 64388 390612 64394
rect 390560 64330 390612 64336
rect 389192 16546 389496 16574
rect 387798 16008 387854 16017
rect 387798 15943 387854 15952
rect 384304 14680 384356 14686
rect 384304 14622 384356 14628
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14622
rect 386696 14612 386748 14618
rect 386696 14554 386748 14560
rect 385960 7676 386012 7682
rect 385960 7618 386012 7624
rect 385972 480 386000 7618
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 14554
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 15943
rect 389468 480 389496 16546
rect 390572 3398 390600 64330
rect 396080 60104 396132 60110
rect 396080 60046 396132 60052
rect 390652 35284 390704 35290
rect 390652 35226 390704 35232
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 35226
rect 391940 29912 391992 29918
rect 391940 29854 391992 29860
rect 391952 16574 391980 29854
rect 391952 16546 392624 16574
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 395344 16040 395396 16046
rect 395344 15982 395396 15988
rect 394240 6316 394292 6322
rect 394240 6258 394292 6264
rect 394252 480 394280 6258
rect 395356 480 395384 15982
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 60046
rect 398840 26988 398892 26994
rect 398840 26930 398892 26936
rect 397460 23112 397512 23118
rect 397460 23054 397512 23060
rect 397472 16574 397500 23054
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3398 398880 26930
rect 402992 16574 403020 75375
rect 408500 71392 408552 71398
rect 408500 71334 408552 71340
rect 407118 20360 407174 20369
rect 407118 20295 407174 20304
rect 404360 18828 404412 18834
rect 404360 18770 404412 18776
rect 402992 16546 403664 16574
rect 398932 15972 398984 15978
rect 398932 15914 398984 15920
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 15914
rect 402520 15904 402572 15910
rect 402520 15846 402572 15852
rect 400864 12096 400916 12102
rect 400864 12038 400916 12044
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 12038
rect 402532 480 402560 15846
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 18770
rect 405738 17368 405794 17377
rect 405738 17303 405794 17312
rect 405752 16574 405780 17303
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3398 407160 20295
rect 408512 16574 408540 71334
rect 412640 67040 412692 67046
rect 412640 66982 412692 66988
rect 409880 29844 409932 29850
rect 409880 29786 409932 29792
rect 409892 16574 409920 29786
rect 411260 27056 411312 27062
rect 411260 26998 411312 27004
rect 411272 16574 411300 26998
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 411272 16546 411944 16574
rect 407210 8936 407266 8945
rect 407210 8871 407266 8880
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 8871
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 66982
rect 415400 61396 415452 61402
rect 415400 61338 415452 61344
rect 414020 25832 414072 25838
rect 414020 25774 414072 25780
rect 414032 16574 414060 25774
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3210 415440 61338
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 415504 3398 415532 57190
rect 425060 50380 425112 50386
rect 425060 50322 425112 50328
rect 418160 49088 418212 49094
rect 418160 49030 418212 49036
rect 416780 29776 416832 29782
rect 416780 29718 416832 29724
rect 416792 16574 416820 29718
rect 418172 16574 418200 49030
rect 422298 29608 422354 29617
rect 422298 29543 422354 29552
rect 419540 17536 419592 17542
rect 419540 17478 419592 17484
rect 419552 16574 419580 17478
rect 422312 16574 422340 29543
rect 423678 17232 423734 17241
rect 423678 17167 423734 17176
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 415412 3182 415532 3210
rect 415504 480 415532 3182
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420918 10296 420974 10305
rect 420918 10231 420974 10240
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 10231
rect 422588 480 422616 16546
rect 423692 3210 423720 17167
rect 425072 16574 425100 50322
rect 426452 16574 426480 80038
rect 430580 79008 430632 79014
rect 430580 78950 430632 78956
rect 427820 60036 427872 60042
rect 427820 59978 427872 59984
rect 427832 16574 427860 59978
rect 430592 16574 430620 78950
rect 462332 78713 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 141642 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 522304 470620 522356 470626
rect 522304 470562 522356 470568
rect 504364 271924 504416 271930
rect 504364 271866 504416 271872
rect 494060 141636 494112 141642
rect 494060 141578 494112 141584
rect 504376 78946 504404 271866
rect 522316 95198 522344 470562
rect 522304 95192 522356 95198
rect 522304 95134 522356 95140
rect 527192 79422 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 558932 141574 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580078 524512 580134 524521
rect 580078 524447 580080 524456
rect 580132 524447 580134 524456
rect 580080 524418 580132 524424
rect 580078 471472 580134 471481
rect 580078 471407 580134 471416
rect 580092 470626 580120 471407
rect 580080 470620 580132 470626
rect 580080 470562 580132 470568
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580092 418198 580120 418231
rect 580080 418192 580132 418198
rect 580080 418134 580132 418140
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580092 378214 580120 378383
rect 580080 378208 580132 378214
rect 580080 378150 580132 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 579986 298752 580042 298761
rect 579986 298687 580042 298696
rect 580000 298178 580028 298687
rect 579988 298172 580040 298178
rect 579988 298114 580040 298120
rect 579986 272232 580042 272241
rect 579986 272167 580042 272176
rect 580000 271930 580028 272167
rect 579988 271924 580040 271930
rect 579988 271866 580040 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 579802 192536 579858 192545
rect 579802 192471 579858 192480
rect 579816 191894 579844 192471
rect 579804 191888 579856 191894
rect 579804 191830 579856 191836
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580000 178090 580028 179143
rect 579988 178084 580040 178090
rect 579988 178026 580040 178032
rect 558920 141568 558972 141574
rect 558920 141510 558972 141516
rect 527180 79416 527232 79422
rect 527180 79358 527232 79364
rect 580092 79354 580120 325207
rect 580184 228410 580212 537775
rect 580172 228404 580224 228410
rect 580172 228346 580224 228352
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 151842 580212 152623
rect 580172 151836 580224 151842
rect 580172 151778 580224 151784
rect 580276 141506 580304 670647
rect 580354 617536 580410 617545
rect 580354 617471 580410 617480
rect 580264 141500 580316 141506
rect 580264 141442 580316 141448
rect 580368 141438 580396 617471
rect 580722 591016 580778 591025
rect 580722 590951 580778 590960
rect 580446 564360 580502 564369
rect 580446 564295 580502 564304
rect 580356 141432 580408 141438
rect 580356 141374 580408 141380
rect 580460 140049 580488 564295
rect 580630 511320 580686 511329
rect 580630 511255 580686 511264
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580446 140040 580502 140049
rect 580446 139975 580502 139984
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580184 125662 580212 125967
rect 580172 125656 580224 125662
rect 580172 125598 580224 125604
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 580552 80714 580580 484599
rect 580644 140146 580672 511255
rect 580736 227050 580764 590951
rect 580906 458144 580962 458153
rect 580906 458079 580962 458088
rect 580814 431624 580870 431633
rect 580814 431559 580870 431568
rect 580724 227044 580776 227050
rect 580724 226986 580776 226992
rect 580632 140140 580684 140146
rect 580632 140082 580684 140088
rect 580540 80708 580592 80714
rect 580540 80650 580592 80656
rect 580828 79393 580856 431559
rect 580920 140078 580948 458079
rect 580908 140072 580960 140078
rect 580908 140014 580960 140020
rect 580814 79384 580870 79393
rect 580080 79348 580132 79354
rect 580814 79319 580870 79328
rect 580080 79290 580132 79296
rect 504364 78940 504416 78946
rect 504364 78882 504416 78888
rect 532700 78872 532752 78878
rect 532700 78814 532752 78820
rect 462318 78704 462374 78713
rect 462318 78639 462374 78648
rect 498200 78124 498252 78130
rect 498200 78066 498252 78072
rect 436742 78024 436798 78033
rect 436742 77959 436798 77968
rect 431960 75472 432012 75478
rect 431960 75414 432012 75420
rect 431972 16574 432000 75414
rect 434720 29708 434772 29714
rect 434720 29650 434772 29656
rect 433340 18760 433392 18766
rect 433340 18702 433392 18708
rect 433352 16574 433380 18702
rect 434732 16574 434760 29650
rect 436100 21548 436152 21554
rect 436100 21490 436152 21496
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 423770 11928 423826 11937
rect 423770 11863 423826 11872
rect 423784 3398 423812 11863
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 7608 429712 7614
rect 429660 7550 429712 7556
rect 429672 480 429700 7550
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 433248 4956 433300 4962
rect 433248 4898 433300 4904
rect 433260 480 433288 4898
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436112 6914 436140 21490
rect 436756 16574 436784 77959
rect 483018 77888 483074 77897
rect 483018 77823 483074 77832
rect 459558 76800 459614 76809
rect 459558 76735 459614 76744
rect 444380 76628 444432 76634
rect 444380 76570 444432 76576
rect 438860 75404 438912 75410
rect 438860 75346 438912 75352
rect 438872 16574 438900 75346
rect 440240 58676 440292 58682
rect 440240 58618 440292 58624
rect 436756 16546 436876 16574
rect 438872 16546 439176 16574
rect 436112 6886 436784 6914
rect 436756 480 436784 6886
rect 436848 5030 436876 16546
rect 436836 5024 436888 5030
rect 436836 4966 436888 4972
rect 437940 3596 437992 3602
rect 437940 3538 437992 3544
rect 437952 480 437980 3538
rect 439148 480 439176 16546
rect 440252 3602 440280 58618
rect 440332 21616 440384 21622
rect 440332 21558 440384 21564
rect 440240 3596 440292 3602
rect 440240 3538 440292 3544
rect 440344 480 440372 21558
rect 442998 21312 443054 21321
rect 442998 21247 443054 21256
rect 441620 17468 441672 17474
rect 441620 17410 441672 17416
rect 441632 16574 441660 17410
rect 443012 16574 443040 21247
rect 444392 16574 444420 76570
rect 447140 35216 447192 35222
rect 447140 35158 447192 35164
rect 445760 20392 445812 20398
rect 445760 20334 445812 20340
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 3596 441580 3602
rect 441528 3538 441580 3544
rect 441540 480 441568 3538
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 20334
rect 447152 16574 447180 35158
rect 454040 28280 454092 28286
rect 454040 28222 454092 28228
rect 449900 20460 449952 20466
rect 449900 20402 449952 20408
rect 448520 20324 448572 20330
rect 448520 20266 448572 20272
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 3482 448560 20266
rect 448612 20256 448664 20262
rect 448612 20198 448664 20204
rect 448624 3602 448652 20198
rect 449912 16574 449940 20402
rect 451280 20188 451332 20194
rect 451280 20130 451332 20136
rect 451292 16574 451320 20130
rect 452660 20120 452712 20126
rect 452660 20062 452712 20068
rect 452672 16574 452700 20062
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3596 448664 3602
rect 448612 3538 448664 3544
rect 449808 3596 449860 3602
rect 449808 3538 449860 3544
rect 448532 3454 448652 3482
rect 448624 480 448652 3454
rect 449820 480 449848 3538
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 28222
rect 456892 20528 456944 20534
rect 456892 20470 456944 20476
rect 456798 20224 456854 20233
rect 456798 20159 456854 20168
rect 455420 20052 455472 20058
rect 455420 19994 455472 20000
rect 455432 16574 455460 19994
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3482 456840 20159
rect 456904 3602 456932 20470
rect 458178 20088 458234 20097
rect 458178 20023 458234 20032
rect 458192 16574 458220 20023
rect 459572 16574 459600 76735
rect 481640 75336 481692 75342
rect 481640 75278 481692 75284
rect 463700 64320 463752 64326
rect 463700 64262 463752 64268
rect 463712 16574 463740 64262
rect 465080 62892 465132 62898
rect 465080 62834 465132 62840
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 456892 3596 456944 3602
rect 456892 3538 456944 3544
rect 458088 3596 458140 3602
rect 458088 3538 458140 3544
rect 456812 3454 456932 3482
rect 456904 480 456932 3454
rect 458100 480 458128 3538
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 462780 3528 462832 3534
rect 461582 3496 461638 3505
rect 462780 3470 462832 3476
rect 461582 3431 461638 3440
rect 461596 480 461624 3431
rect 462792 480 462820 3470
rect 463988 480 464016 16546
rect 465092 3534 465120 62834
rect 474002 35184 474058 35193
rect 474002 35119 474058 35128
rect 466460 32428 466512 32434
rect 466460 32370 466512 32376
rect 465172 31204 465224 31210
rect 465172 31146 465224 31152
rect 465080 3528 465132 3534
rect 465080 3470 465132 3476
rect 465184 480 465212 31146
rect 466472 16574 466500 32370
rect 467840 23044 467892 23050
rect 467840 22986 467892 22992
rect 467852 16574 467880 22986
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 465908 3528 465960 3534
rect 465908 3470 465960 3476
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465920 354 465948 3470
rect 467484 480 467512 16546
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 473358 15872 473414 15881
rect 473358 15807 473414 15816
rect 469864 10396 469916 10402
rect 469864 10338 469916 10344
rect 469876 480 469904 10338
rect 471060 6248 471112 6254
rect 471060 6190 471112 6196
rect 471072 480 471100 6190
rect 473372 3534 473400 15807
rect 473452 12028 473504 12034
rect 473452 11970 473504 11976
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 472254 3360 472310 3369
rect 472254 3295 472310 3304
rect 472268 480 472296 3295
rect 473464 480 473492 11970
rect 474016 3602 474044 35119
rect 477498 22808 477554 22817
rect 477498 22743 477554 22752
rect 476118 19952 476174 19961
rect 476118 19887 476174 19896
rect 476132 16574 476160 19887
rect 477512 16574 477540 22743
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 474004 3596 474056 3602
rect 474004 3538 474056 3544
rect 474188 3528 474240 3534
rect 474188 3470 474240 3476
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3470
rect 475752 3460 475804 3466
rect 475752 3402 475804 3408
rect 475764 480 475792 3402
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 4956 479392 4962
rect 479340 4898 479392 4904
rect 479352 480 479380 4898
rect 480536 4888 480588 4894
rect 480536 4830 480588 4836
rect 480548 480 480576 4830
rect 481652 3466 481680 75278
rect 481732 19984 481784 19990
rect 481732 19926 481784 19932
rect 481640 3460 481692 3466
rect 481640 3402 481692 3408
rect 481744 480 481772 19926
rect 483032 16574 483060 77823
rect 496818 75304 496874 75313
rect 489920 75268 489972 75274
rect 496818 75239 496874 75248
rect 489920 75210 489972 75216
rect 487160 64252 487212 64258
rect 487160 64194 487212 64200
rect 485780 49020 485832 49026
rect 485780 48962 485832 48968
rect 484400 21480 484452 21486
rect 484400 21422 484452 21428
rect 484412 16574 484440 21422
rect 485792 16574 485820 48962
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 482468 3460 482520 3466
rect 482468 3402 482520 3408
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3402
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 64194
rect 488816 13116 488868 13122
rect 488816 13058 488868 13064
rect 488828 480 488856 13058
rect 489932 480 489960 75210
rect 490012 71324 490064 71330
rect 490012 71266 490064 71272
rect 490024 16574 490052 71266
rect 491300 21412 491352 21418
rect 491300 21354 491352 21360
rect 491312 16574 491340 21354
rect 492680 17400 492732 17406
rect 492680 17342 492732 17348
rect 492692 16574 492720 17342
rect 496832 16574 496860 75239
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494702 5128 494758 5137
rect 494702 5063 494758 5072
rect 494716 480 494744 5063
rect 495900 3528 495952 3534
rect 495900 3470 495952 3476
rect 495912 480 495940 3470
rect 497108 480 497136 16546
rect 498212 480 498240 78066
rect 505098 76664 505154 76673
rect 505098 76599 505154 76608
rect 500958 72448 501014 72457
rect 500958 72383 501014 72392
rect 500972 16574 501000 72383
rect 503720 17332 503772 17338
rect 503720 17274 503772 17280
rect 500972 16546 501368 16574
rect 500592 14544 500644 14550
rect 500592 14486 500644 14492
rect 498936 11960 498988 11966
rect 498936 11902 498988 11908
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 11902
rect 500604 480 500632 14486
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502984 11892 503036 11898
rect 502984 11834 503036 11840
rect 502996 480 503024 11834
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 17274
rect 505112 16574 505140 76599
rect 507860 71256 507912 71262
rect 507860 71198 507912 71204
rect 507872 16574 507900 71198
rect 523040 71188 523092 71194
rect 523040 71130 523092 71136
rect 518900 69760 518952 69766
rect 518900 69702 518952 69708
rect 514760 62824 514812 62830
rect 514760 62766 514812 62772
rect 511998 55856 512054 55865
rect 511998 55791 512054 55800
rect 505112 16546 505416 16574
rect 507872 16546 508912 16574
rect 505388 480 505416 16546
rect 506480 11824 506532 11830
rect 506480 11766 506532 11772
rect 506492 480 506520 11766
rect 507676 9036 507728 9042
rect 507676 8978 507728 8984
rect 507688 480 507716 8978
rect 508884 480 508912 16546
rect 511262 14512 511318 14521
rect 511262 14447 511318 14456
rect 509608 11756 509660 11762
rect 509608 11698 509660 11704
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 11698
rect 511276 480 511304 14447
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 55791
rect 513378 11792 513434 11801
rect 513378 11727 513434 11736
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 11727
rect 514772 3534 514800 62766
rect 516140 22976 516192 22982
rect 516140 22918 516192 22924
rect 514852 17264 514904 17270
rect 514852 17206 514904 17212
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 17206
rect 516152 16574 516180 22918
rect 518912 16574 518940 69702
rect 520280 22908 520332 22914
rect 520280 22850 520332 22856
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 518348 4820 518400 4826
rect 518348 4762 518400 4768
rect 518360 480 518388 4762
rect 519556 480 519584 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 22850
rect 521844 8968 521896 8974
rect 521844 8910 521896 8916
rect 521856 480 521884 8910
rect 523052 480 523080 71130
rect 529938 66872 529994 66881
rect 529938 66807 529994 66816
rect 525800 65612 525852 65618
rect 525800 65554 525852 65560
rect 524420 31136 524472 31142
rect 524420 31078 524472 31084
rect 524432 16574 524460 31078
rect 525812 16574 525840 65554
rect 527180 22840 527232 22846
rect 527180 22782 527232 22788
rect 527192 16574 527220 22782
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523776 14476 523828 14482
rect 523776 14418 523828 14424
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 14418
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 528558 13016 528614 13025
rect 528558 12951 528614 12960
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 12951
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 66807
rect 531318 28248 531374 28257
rect 531318 28183 531374 28192
rect 531332 3534 531360 28183
rect 531410 18728 531466 18737
rect 531410 18663 531466 18672
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 18663
rect 532712 16574 532740 78814
rect 554780 78804 554832 78810
rect 554780 78746 554832 78752
rect 549258 75168 549314 75177
rect 549258 75103 549314 75112
rect 536840 71120 536892 71126
rect 536840 71062 536892 71068
rect 535460 31068 535512 31074
rect 535460 31010 535512 31016
rect 534080 24472 534132 24478
rect 534080 24414 534132 24420
rect 534092 16574 534120 24414
rect 535472 16574 535500 31010
rect 536852 16574 536880 71062
rect 539600 71052 539652 71058
rect 539600 70994 539652 71000
rect 538220 24404 538272 24410
rect 538220 24346 538272 24352
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 24346
rect 539612 3534 539640 70994
rect 543740 66972 543792 66978
rect 543740 66914 543792 66920
rect 542360 29640 542412 29646
rect 542360 29582 542412 29588
rect 540980 24336 541032 24342
rect 540980 24278 541032 24284
rect 540992 16574 541020 24278
rect 542372 16574 542400 29582
rect 543752 16574 543780 66914
rect 545120 24268 545172 24274
rect 545120 24210 545172 24216
rect 545132 16574 545160 24210
rect 546498 18592 546554 18601
rect 546498 18527 546554 18536
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 539692 10328 539744 10334
rect 539692 10270 539744 10276
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 10270
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 18527
rect 549272 16574 549300 75103
rect 550638 42120 550694 42129
rect 550638 42055 550694 42064
rect 550652 16574 550680 42055
rect 552020 24200 552072 24206
rect 552020 24142 552072 24148
rect 552032 16574 552060 24142
rect 553400 18692 553452 18698
rect 553400 18634 553452 18640
rect 553412 16574 553440 18634
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 549074 6352 549130 6361
rect 549074 6287 549130 6296
rect 547878 4992 547934 5001
rect 547878 4927 547934 4936
rect 547892 480 547920 4927
rect 549088 480 549116 6287
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 78746
rect 557540 78736 557592 78742
rect 557540 78678 557592 78684
rect 556160 25764 556212 25770
rect 556160 25706 556212 25712
rect 556172 480 556200 25706
rect 556252 18624 556304 18630
rect 556252 18566 556304 18572
rect 556264 16574 556292 18566
rect 557552 16574 557580 78678
rect 574744 78056 574796 78062
rect 574744 77998 574796 78004
rect 558920 76560 558972 76566
rect 558920 76502 558972 76508
rect 565818 76528 565874 76537
rect 558932 16574 558960 76502
rect 565818 76463 565874 76472
rect 564440 75200 564492 75206
rect 564440 75142 564492 75148
rect 560300 26920 560352 26926
rect 560300 26862 560352 26868
rect 560312 16574 560340 26862
rect 563060 25696 563112 25702
rect 563060 25638 563112 25644
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562048 6180 562100 6186
rect 562048 6122 562100 6128
rect 562060 480 562088 6122
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 25638
rect 564452 480 564480 75142
rect 564532 69692 564584 69698
rect 564532 69634 564584 69640
rect 564544 16574 564572 69634
rect 565832 16574 565860 76463
rect 569960 66904 570012 66910
rect 569960 66846 570012 66852
rect 568580 64184 568632 64190
rect 568580 64126 568632 64132
rect 567198 30968 567254 30977
rect 567198 30903 567254 30912
rect 567212 16574 567240 30903
rect 568592 16574 568620 64126
rect 569972 16574 570000 66846
rect 572720 65544 572772 65550
rect 572720 65486 572772 65492
rect 571340 25628 571392 25634
rect 571340 25570 571392 25576
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 25570
rect 572732 480 572760 65486
rect 572812 25560 572864 25566
rect 572812 25502 572864 25508
rect 572824 16574 572852 25502
rect 572824 16546 573496 16574
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 574650 11656 574706 11665
rect 574650 11591 574706 11600
rect 574664 3482 574692 11591
rect 574756 3602 574784 77998
rect 581092 77988 581144 77994
rect 581092 77930 581144 77936
rect 578238 73808 578294 73817
rect 578238 73743 578294 73752
rect 578252 16574 578280 73743
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579620 24132 579672 24138
rect 579620 24074 579672 24080
rect 579632 19825 579660 24074
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579618 19816 579674 19825
rect 579618 19751 579674 19760
rect 578252 16546 578648 16574
rect 576306 6216 576362 6225
rect 576306 6151 576362 6160
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 576320 480 576348 6151
rect 577410 4856 577466 4865
rect 577410 4791 577466 4800
rect 577424 480 577452 4791
rect 578620 480 578648 16546
rect 580276 6633 580304 22714
rect 581104 16574 581132 77930
rect 582378 22672 582434 22681
rect 582378 22607 582434 22616
rect 582392 16574 582420 22607
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 2778 579964 2834 580000
rect 2778 579944 2780 579964
rect 2780 579944 2832 579964
rect 2832 579944 2834 579964
rect 3054 566888 3110 566944
rect 3330 423544 3386 423600
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3146 319232 3202 319288
rect 3330 306176 3386 306232
rect 3238 293120 3294 293176
rect 3146 267144 3202 267200
rect 3238 254088 3294 254144
rect 3238 241032 3294 241088
rect 3238 227976 3294 228032
rect 3238 214920 3294 214976
rect 3238 201864 3294 201920
rect 3146 188808 3202 188864
rect 3146 162868 3148 162888
rect 3148 162868 3200 162888
rect 3200 162868 3202 162888
rect 3146 162832 3202 162868
rect 3330 149776 3386 149832
rect 3146 110608 3202 110664
rect 3330 136720 3386 136776
rect 3238 97552 3294 97608
rect 3146 84632 3202 84688
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3606 606056 3662 606112
rect 3514 527876 3570 527912
rect 3514 527856 3516 527876
rect 3516 527856 3568 527876
rect 3568 527856 3570 527876
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 475632 3570 475688
rect 3514 462576 3570 462632
rect 3514 449520 3570 449576
rect 3790 553832 3846 553888
rect 3698 397432 3754 397488
rect 3974 501744 4030 501800
rect 3882 345344 3938 345400
rect 4066 358400 4122 358456
rect 6918 79464 6974 79520
rect 3974 79328 4030 79384
rect 3790 79192 3846 79248
rect 3606 79056 3662 79112
rect 3422 78920 3478 78976
rect 2778 75248 2834 75304
rect 1398 75112 1454 75168
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 3330 19352 3386 19408
rect 3422 6432 3478 6488
rect 4066 4800 4122 4856
rect 10322 77832 10378 77888
rect 45006 141344 45062 141400
rect 44914 80416 44970 80472
rect 116674 130056 116730 130112
rect 118238 136040 118294 136096
rect 117318 133320 117374 133376
rect 116950 132232 117006 132288
rect 116858 131144 116914 131200
rect 117318 128968 117374 129024
rect 117318 127880 117374 127936
rect 117686 126792 117742 126848
rect 117318 125704 117374 125760
rect 117870 125704 117926 125760
rect 117778 123528 117834 123584
rect 117686 122440 117742 122496
rect 117410 121352 117466 121408
rect 117318 120264 117374 120320
rect 117870 119176 117926 119232
rect 117318 118088 117374 118144
rect 117318 117000 117374 117056
rect 117410 115912 117466 115968
rect 117318 114824 117374 114880
rect 117318 113736 117374 113792
rect 117318 112648 117374 112704
rect 117318 111560 117374 111616
rect 117410 110472 117466 110528
rect 117318 109384 117374 109440
rect 117318 108296 117374 108352
rect 117318 107208 117374 107264
rect 117318 106120 117374 106176
rect 117410 105032 117466 105088
rect 117318 103944 117374 104000
rect 118054 94152 118110 94208
rect 118146 91976 118202 92032
rect 118422 136604 118478 136640
rect 118422 136584 118424 136604
rect 118424 136584 118476 136604
rect 118476 136584 118478 136604
rect 118422 134952 118478 135008
rect 118330 93064 118386 93120
rect 118238 90888 118294 90944
rect 118422 89800 118478 89856
rect 118606 102856 118662 102912
rect 138110 195916 138112 195936
rect 138112 195916 138164 195936
rect 138164 195916 138166 195936
rect 138110 195880 138166 195916
rect 140410 195880 140466 195936
rect 140778 195608 140834 195664
rect 139398 195472 139454 195528
rect 149610 193296 149666 193352
rect 140778 191800 140834 191856
rect 140962 191664 141018 191720
rect 140870 191528 140926 191584
rect 140778 190848 140834 190904
rect 119158 101768 119214 101824
rect 119250 100680 119306 100736
rect 119066 99592 119122 99648
rect 118974 98504 119030 98560
rect 118882 97416 118938 97472
rect 118790 95240 118846 95296
rect 118698 88712 118754 88768
rect 118514 87624 118570 87680
rect 118514 86536 118570 86592
rect 118238 84360 118294 84416
rect 44822 78512 44878 78568
rect 37278 76608 37334 76664
rect 20718 76472 20774 76528
rect 20626 3304 20682 3360
rect 23018 7520 23074 7576
rect 35898 73752 35954 73808
rect 41878 8880 41934 8936
rect 40682 6160 40738 6216
rect 57978 74024 58034 74080
rect 53838 73888 53894 73944
rect 57242 9152 57298 9208
rect 56046 9016 56102 9072
rect 71778 74160 71834 74216
rect 74998 10240 75054 10296
rect 73802 6296 73858 6352
rect 91098 44784 91154 44840
rect 92478 10376 92534 10432
rect 109314 7656 109370 7712
rect 111798 76744 111854 76800
rect 110510 10512 110566 10568
rect 118330 83272 118386 83328
rect 118606 85448 118662 85504
rect 139398 187584 139454 187640
rect 140778 186224 140834 186280
rect 140778 182552 140834 182608
rect 165434 193296 165490 193352
rect 140962 182688 141018 182744
rect 140870 182416 140926 182472
rect 144642 180920 144698 180976
rect 146022 180956 146024 180976
rect 146024 180956 146076 180976
rect 146076 180956 146078 180976
rect 146022 180920 146078 180956
rect 144090 178880 144146 178936
rect 141606 178744 141662 178800
rect 142066 178608 142122 178664
rect 141698 178472 141754 178528
rect 142526 172896 142582 172952
rect 149334 175344 149390 175400
rect 154394 175380 154396 175400
rect 154396 175380 154448 175400
rect 154448 175380 154450 175400
rect 154394 175344 154450 175380
rect 155222 156576 155278 156632
rect 165434 175480 165490 175536
rect 171138 174528 171194 174584
rect 165434 172896 165490 172952
rect 120630 136040 120686 136096
rect 120538 134952 120594 135008
rect 119342 77968 119398 78024
rect 179510 128152 179566 128208
rect 179418 126792 179474 126848
rect 125230 80144 125286 80200
rect 124770 79872 124826 79928
rect 122102 78104 122158 78160
rect 123666 75248 123722 75304
rect 125046 77832 125102 77888
rect 125322 79736 125378 79792
rect 126104 79872 126160 79928
rect 126564 79872 126620 79928
rect 126748 79906 126804 79962
rect 125506 77832 125562 77888
rect 125598 75112 125654 75168
rect 125782 77696 125838 77752
rect 127116 79906 127172 79962
rect 127300 79906 127356 79962
rect 127576 79872 127632 79928
rect 127760 79906 127816 79962
rect 127162 76472 127218 76528
rect 127346 78104 127402 78160
rect 128312 79872 128368 79928
rect 128680 79872 128736 79928
rect 129232 79872 129288 79928
rect 127438 77832 127494 77888
rect 127990 79600 128046 79656
rect 128266 79600 128322 79656
rect 128726 79636 128728 79656
rect 128728 79636 128780 79656
rect 128780 79636 128782 79656
rect 128358 78784 128414 78840
rect 128726 79600 128782 79636
rect 128450 76608 128506 76664
rect 129876 79872 129932 79928
rect 130060 79872 130116 79928
rect 129370 78648 129426 78704
rect 129738 78784 129794 78840
rect 129738 77832 129794 77888
rect 130014 78648 130070 78704
rect 131164 79906 131220 79962
rect 131348 79872 131404 79928
rect 130382 74432 130438 74488
rect 131210 78648 131266 78704
rect 131670 78104 131726 78160
rect 132176 79906 132232 79962
rect 132544 79906 132600 79962
rect 132774 79736 132830 79792
rect 133004 79906 133060 79962
rect 132682 79636 132684 79656
rect 132684 79636 132736 79656
rect 132736 79636 132738 79656
rect 132682 79600 132738 79636
rect 132590 77968 132646 78024
rect 133924 79872 133980 79928
rect 134292 79872 134348 79928
rect 134476 79906 134532 79962
rect 134430 79736 134486 79792
rect 134752 79872 134808 79928
rect 134936 79906 134992 79962
rect 134338 79600 134394 79656
rect 134062 78648 134118 78704
rect 133970 77968 134026 78024
rect 134338 76744 134394 76800
rect 134798 79600 134854 79656
rect 134982 79736 135038 79792
rect 135396 79872 135452 79928
rect 135672 79872 135728 79928
rect 136500 79906 136556 79962
rect 136776 79906 136832 79962
rect 135810 79600 135866 79656
rect 136454 79736 136510 79792
rect 136960 79906 137016 79962
rect 136638 79600 136694 79656
rect 136822 78784 136878 78840
rect 137006 79736 137062 79792
rect 137236 79872 137292 79928
rect 137420 79906 137476 79962
rect 138064 79872 138120 79928
rect 137926 79736 137982 79792
rect 137374 79600 137430 79656
rect 137926 79600 137982 79656
rect 138110 78784 138166 78840
rect 138018 78648 138074 78704
rect 139076 79906 139132 79962
rect 139030 79600 139086 79656
rect 139444 79906 139500 79962
rect 140088 79838 140144 79894
rect 139352 79770 139408 79826
rect 139950 79736 140006 79792
rect 139122 78648 139178 78704
rect 139582 79600 139638 79656
rect 139398 75928 139454 75984
rect 140042 79600 140098 79656
rect 140916 79906 140972 79962
rect 141284 79872 141340 79928
rect 141560 79906 141616 79962
rect 141928 79872 141984 79928
rect 142112 79906 142168 79962
rect 140594 75792 140650 75848
rect 140962 79600 141018 79656
rect 140870 78784 140926 78840
rect 140686 75520 140742 75576
rect 140502 73072 140558 73128
rect 141422 79600 141478 79656
rect 141606 79736 141662 79792
rect 141606 78104 141662 78160
rect 141974 79736 142030 79792
rect 141790 76336 141846 76392
rect 142480 79838 142536 79894
rect 142342 79600 142398 79656
rect 141974 77016 142030 77072
rect 142940 79906 142996 79962
rect 143400 79872 143456 79928
rect 143308 79736 143364 79792
rect 144136 79906 144192 79962
rect 142894 77696 142950 77752
rect 142434 3984 142490 4040
rect 142342 3848 142398 3904
rect 143262 76608 143318 76664
rect 144504 79872 144560 79928
rect 144688 79906 144744 79962
rect 145516 79872 145572 79928
rect 143446 74024 143502 74080
rect 143814 79600 143870 79656
rect 143814 77152 143870 77208
rect 143814 76608 143870 76664
rect 144458 79600 144514 79656
rect 144550 77832 144606 77888
rect 145332 79736 145388 79792
rect 145286 79600 145342 79656
rect 144918 75928 144974 75984
rect 144642 73888 144698 73944
rect 143078 3168 143134 3224
rect 146068 79872 146124 79928
rect 145746 79620 145802 79656
rect 145746 79600 145748 79620
rect 145748 79600 145800 79620
rect 145800 79600 145802 79620
rect 146344 79906 146400 79962
rect 146528 79838 146584 79894
rect 147356 79906 147412 79962
rect 147540 79906 147596 79962
rect 147310 79772 147312 79792
rect 147312 79772 147364 79792
rect 147364 79772 147366 79792
rect 147310 79736 147366 79772
rect 147586 79736 147642 79792
rect 147816 79906 147872 79962
rect 146022 75792 146078 75848
rect 146298 79600 146354 79656
rect 146206 74160 146262 74216
rect 144550 3440 144606 3496
rect 147126 79600 147182 79656
rect 147310 76200 147366 76256
rect 147862 79736 147918 79792
rect 147770 79600 147826 79656
rect 147586 77152 147642 77208
rect 147494 75928 147550 75984
rect 148368 79872 148424 79928
rect 148046 76608 148102 76664
rect 148552 79906 148608 79962
rect 148828 79906 148884 79962
rect 149012 79736 149068 79792
rect 149472 79906 149528 79962
rect 150300 79906 150356 79962
rect 148690 76744 148746 76800
rect 148966 79600 149022 79656
rect 148782 76608 148838 76664
rect 150208 79736 150264 79792
rect 149978 78104 150034 78160
rect 150852 79872 150908 79928
rect 150070 77288 150126 77344
rect 150530 78104 150586 78160
rect 151496 79906 151552 79962
rect 151358 79736 151414 79792
rect 151680 79736 151736 79792
rect 151864 79872 151920 79928
rect 151726 78784 151782 78840
rect 151542 78648 151598 78704
rect 151910 78648 151966 78704
rect 152600 79872 152656 79928
rect 152876 79906 152932 79962
rect 152922 79736 152978 79792
rect 153152 79906 153208 79962
rect 153106 79600 153162 79656
rect 152922 77288 152978 77344
rect 146850 3984 146906 4040
rect 146850 3576 146906 3632
rect 153934 79736 153990 79792
rect 154532 79872 154588 79928
rect 154486 79736 154542 79792
rect 154394 79600 154450 79656
rect 155728 79872 155784 79928
rect 156188 79906 156244 79962
rect 156372 79906 156428 79962
rect 157108 79906 157164 79962
rect 157292 79906 157348 79962
rect 155958 79600 156014 79656
rect 155866 76880 155922 76936
rect 156234 75248 156290 75304
rect 156602 79600 156658 79656
rect 156694 75112 156750 75168
rect 156970 78648 157026 78704
rect 157568 79736 157624 79792
rect 157798 79736 157854 79792
rect 158120 79872 158176 79928
rect 158304 79872 158360 79928
rect 158580 79906 158636 79962
rect 158948 79838 159004 79894
rect 159316 79872 159372 79928
rect 159500 79872 159556 79928
rect 157154 75384 157210 75440
rect 157890 79620 157946 79656
rect 157890 79600 157892 79620
rect 157892 79600 157944 79620
rect 157944 79600 157946 79620
rect 157798 77288 157854 77344
rect 158718 79600 158774 79656
rect 158442 76608 158498 76664
rect 158350 74432 158406 74488
rect 159270 79600 159326 79656
rect 159178 77832 159234 77888
rect 159454 79600 159510 79656
rect 159776 79906 159832 79962
rect 160236 79872 160292 79928
rect 159822 79736 159878 79792
rect 160098 79600 160154 79656
rect 160282 78784 160338 78840
rect 160190 75928 160246 75984
rect 160374 75928 160430 75984
rect 160880 79872 160936 79928
rect 161064 79872 161120 79928
rect 161432 79906 161488 79962
rect 161616 79872 161672 79928
rect 160926 79772 160928 79792
rect 160928 79772 160980 79792
rect 160980 79772 160982 79792
rect 160926 79736 160982 79772
rect 161110 79636 161112 79656
rect 161112 79636 161164 79656
rect 161164 79636 161166 79656
rect 160742 78648 160798 78704
rect 161110 79600 161166 79636
rect 160650 75792 160706 75848
rect 161294 78104 161350 78160
rect 161386 76744 161442 76800
rect 160098 6160 160154 6216
rect 158902 4800 158958 4856
rect 162444 79824 162500 79826
rect 162444 79772 162446 79824
rect 162446 79772 162498 79824
rect 162498 79772 162500 79824
rect 162444 79770 162500 79772
rect 162674 79636 162676 79656
rect 162676 79636 162728 79656
rect 162728 79636 162730 79656
rect 162030 75792 162086 75848
rect 162674 79600 162730 79636
rect 162398 75792 162454 75848
rect 162674 77832 162730 77888
rect 162858 79736 162914 79792
rect 162950 78240 163006 78296
rect 162858 76200 162914 76256
rect 162766 75928 162822 75984
rect 163732 79872 163788 79928
rect 164100 79906 164156 79962
rect 163686 79736 163742 79792
rect 163502 79600 163558 79656
rect 163410 78648 163466 78704
rect 164054 79636 164056 79656
rect 164056 79636 164108 79656
rect 164108 79636 164110 79656
rect 164054 79600 164110 79636
rect 164560 79906 164616 79962
rect 164744 79906 164800 79962
rect 165020 79906 165076 79962
rect 164146 75248 164202 75304
rect 164790 79600 164846 79656
rect 165480 79872 165536 79928
rect 166032 79872 166088 79928
rect 166216 79872 166272 79928
rect 165066 79600 165122 79656
rect 165158 76608 165214 76664
rect 165342 75928 165398 75984
rect 165526 78784 165582 78840
rect 165618 77288 165674 77344
rect 165986 75928 166042 75984
rect 166952 79872 167008 79928
rect 166538 75928 166594 75984
rect 166906 79600 166962 79656
rect 167320 79906 167376 79962
rect 168240 79872 168296 79928
rect 166722 73208 166778 73264
rect 166906 76064 166962 76120
rect 168010 79736 168066 79792
rect 168378 79772 168380 79792
rect 168380 79772 168432 79792
rect 168432 79772 168434 79792
rect 168102 79464 168158 79520
rect 168102 78648 168158 78704
rect 168194 77424 168250 77480
rect 168010 75928 168066 75984
rect 168378 79736 168434 79772
rect 168286 75112 168342 75168
rect 168792 79906 168848 79962
rect 168976 79906 169032 79962
rect 169896 79872 169952 79928
rect 168746 79600 168802 79656
rect 169436 79736 169492 79792
rect 169850 79736 169906 79792
rect 170448 79906 170504 79962
rect 169390 79600 169446 79656
rect 169666 79600 169722 79656
rect 169666 76472 169722 76528
rect 169942 77424 169998 77480
rect 170816 79736 170872 79792
rect 171092 79872 171148 79928
rect 171368 79906 171424 79962
rect 170494 77424 170550 77480
rect 170402 77288 170458 77344
rect 169758 11600 169814 11656
rect 171138 79600 171194 79656
rect 171552 79872 171608 79928
rect 171138 78240 171194 78296
rect 171138 77968 171194 78024
rect 171506 78920 171562 78976
rect 172196 79906 172252 79962
rect 172380 79872 172436 79928
rect 171782 79056 171838 79112
rect 171782 78240 171838 78296
rect 173024 79872 173080 79928
rect 173300 79906 173356 79962
rect 172978 79756 173034 79792
rect 172978 79736 172980 79756
rect 172980 79736 173032 79756
rect 173032 79736 173034 79756
rect 172518 79464 172574 79520
rect 172242 78920 172298 78976
rect 171690 77696 171746 77752
rect 172702 78784 172758 78840
rect 173944 79872 174000 79928
rect 173990 79736 174046 79792
rect 173162 78240 173218 78296
rect 173530 79328 173586 79384
rect 173714 78920 173770 78976
rect 173162 76336 173218 76392
rect 172518 61376 172574 61432
rect 173254 69536 173310 69592
rect 173898 75656 173954 75712
rect 174358 79600 174414 79656
rect 176290 79328 176346 79384
rect 176106 79056 176162 79112
rect 175922 78784 175978 78840
rect 175646 78648 175702 78704
rect 180890 129648 180946 129704
rect 180798 125568 180854 125624
rect 180430 79464 180486 79520
rect 174542 77696 174598 77752
rect 176658 62736 176714 62792
rect 180062 75792 180118 75848
rect 181074 131008 181130 131064
rect 180982 107888 181038 107944
rect 182178 124208 182234 124264
rect 182730 120128 182786 120184
rect 182638 118768 182694 118824
rect 182546 117408 182602 117464
rect 182454 116048 182510 116104
rect 182362 114688 182418 114744
rect 182270 113328 182326 113384
rect 183006 122848 183062 122904
rect 182914 121488 182970 121544
rect 182822 111968 182878 112024
rect 182178 109248 182234 109304
rect 182270 88848 182326 88904
rect 183282 106528 183338 106584
rect 183282 105168 183338 105224
rect 183282 103808 183338 103864
rect 183282 102448 183338 102504
rect 183282 101088 183338 101144
rect 183190 99728 183246 99784
rect 183190 98368 183246 98424
rect 183190 97008 183246 97064
rect 183190 95648 183246 95704
rect 183466 94288 183522 94344
rect 183466 92928 183522 92984
rect 183466 91568 183522 91624
rect 183466 90208 183522 90264
rect 182822 87488 182878 87544
rect 182730 86128 182786 86184
rect 182730 84768 182786 84824
rect 182730 83408 182786 83464
rect 182914 82048 182970 82104
rect 182822 80688 182878 80744
rect 393962 80552 394018 80608
rect 194598 75520 194654 75576
rect 193218 65456 193274 65512
rect 191838 17040 191894 17096
rect 194414 6024 194470 6080
rect 197910 8744 197966 8800
rect 212538 34040 212594 34096
rect 210974 3984 211030 4040
rect 214470 3168 214526 3224
rect 218150 3848 218206 3904
rect 221554 3712 221610 3768
rect 230478 74024 230534 74080
rect 226430 33904 226486 33960
rect 229374 13232 229430 13288
rect 228730 6840 228786 6896
rect 255962 78104 256018 78160
rect 244278 73888 244334 73944
rect 242898 26968 242954 27024
rect 235814 3576 235870 3632
rect 248418 20440 248474 20496
rect 246394 6704 246450 6760
rect 282918 77152 282974 77208
rect 251178 17856 251234 17912
rect 266358 33768 266414 33824
rect 280158 17720 280214 17776
rect 264978 14864 265034 14920
rect 264150 6568 264206 6624
rect 279054 14728 279110 14784
rect 281906 9560 281962 9616
rect 284390 17584 284446 17640
rect 298098 72528 298154 72584
rect 300858 17448 300914 17504
rect 354678 77016 354734 77072
rect 299662 9424 299718 9480
rect 300766 6432 300822 6488
rect 316038 35264 316094 35320
rect 317418 26832 317474 26888
rect 315026 9288 315082 9344
rect 317326 9152 317382 9208
rect 336738 31048 336794 31104
rect 335358 28328 335414 28384
rect 334622 12008 334678 12064
rect 353298 68176 353354 68232
rect 351918 51720 351974 51776
rect 351642 9016 351698 9072
rect 372618 58520 372674 58576
rect 365718 16088 365774 16144
rect 370134 14592 370190 14648
rect 371238 13096 371294 13152
rect 397458 78784 397514 78840
rect 389178 76880 389234 76936
rect 402978 75384 403034 75440
rect 387798 15952 387854 16008
rect 407118 20304 407174 20360
rect 405738 17312 405794 17368
rect 407210 8880 407266 8936
rect 422298 29552 422354 29608
rect 423678 17176 423734 17232
rect 420918 10240 420974 10296
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 577632 580226 577688
rect 580170 537784 580226 537840
rect 580078 524476 580134 524512
rect 580078 524456 580080 524476
rect 580080 524456 580132 524476
rect 580132 524456 580134 524476
rect 580078 471416 580134 471472
rect 580078 418240 580134 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 579802 365064 579858 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 325216 580134 325272
rect 579986 312024 580042 312080
rect 579986 298696 580042 298752
rect 579986 272176 580042 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 579802 232328 579858 232384
rect 579802 192480 579858 192536
rect 579986 179152 580042 179208
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580354 617480 580410 617536
rect 580722 590960 580778 591016
rect 580446 564304 580502 564360
rect 580630 511264 580686 511320
rect 580538 484608 580594 484664
rect 580446 139984 580502 140040
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580906 458088 580962 458144
rect 580814 431568 580870 431624
rect 580814 79328 580870 79384
rect 462318 78648 462374 78704
rect 436742 77968 436798 78024
rect 423770 11872 423826 11928
rect 483018 77832 483074 77888
rect 459558 76744 459614 76800
rect 442998 21256 443054 21312
rect 456798 20168 456854 20224
rect 458178 20032 458234 20088
rect 461582 3440 461638 3496
rect 474002 35128 474058 35184
rect 473358 15816 473414 15872
rect 472254 3304 472310 3360
rect 477498 22752 477554 22808
rect 476118 19896 476174 19952
rect 496818 75248 496874 75304
rect 494702 5072 494758 5128
rect 505098 76608 505154 76664
rect 500958 72392 501014 72448
rect 511998 55800 512054 55856
rect 511262 14456 511318 14512
rect 513378 11736 513434 11792
rect 529938 66816 529994 66872
rect 528558 12960 528614 13016
rect 531318 28192 531374 28248
rect 531410 18672 531466 18728
rect 549258 75112 549314 75168
rect 546498 18536 546554 18592
rect 550638 42064 550694 42120
rect 549074 6296 549130 6352
rect 547878 4936 547934 4992
rect 565818 76472 565874 76528
rect 567198 30912 567254 30968
rect 574650 11600 574706 11656
rect 578238 73752 578294 73808
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579618 19760 579674 19816
rect 576306 6160 576362 6216
rect 577410 4800 577466 4856
rect 582378 22616 582434 22672
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580349 617538 580415 617541
rect 583520 617538 584960 617628
rect 580349 617536 584960 617538
rect 580349 617480 580354 617536
rect 580410 617480 584960 617536
rect 580349 617478 584960 617480
rect 580349 617475 580415 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580717 591018 580783 591021
rect 583520 591018 584960 591108
rect 580717 591016 584960 591018
rect 580717 590960 580722 591016
rect 580778 590960 584960 591016
rect 580717 590958 584960 590960
rect 580717 590955 580783 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 2773 580002 2839 580005
rect -960 580000 2839 580002
rect -960 579944 2778 580000
rect 2834 579944 2839 580000
rect -960 579942 2839 579944
rect -960 579852 480 579942
rect 2773 579939 2839 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580441 564362 580507 564365
rect 583520 564362 584960 564452
rect 580441 564360 584960 564362
rect 580441 564304 580446 564360
rect 580502 564304 584960 564360
rect 580441 564302 584960 564304
rect 580441 564299 580507 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3785 553890 3851 553893
rect -960 553888 3851 553890
rect -960 553832 3790 553888
rect 3846 553832 3851 553888
rect -960 553830 3851 553832
rect -960 553740 480 553830
rect 3785 553827 3851 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 580073 524514 580139 524517
rect 583520 524514 584960 524604
rect 580073 524512 584960 524514
rect 580073 524456 580078 524512
rect 580134 524456 584960 524512
rect 580073 524454 584960 524456
rect 580073 524451 580139 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580625 511322 580691 511325
rect 583520 511322 584960 511412
rect 580625 511320 584960 511322
rect 580625 511264 580630 511320
rect 580686 511264 584960 511320
rect 580625 511262 584960 511264
rect 580625 511259 580691 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3969 501802 4035 501805
rect -960 501800 4035 501802
rect -960 501744 3974 501800
rect 4030 501744 4035 501800
rect -960 501742 4035 501744
rect -960 501652 480 501742
rect 3969 501739 4035 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 580073 471474 580139 471477
rect 583520 471474 584960 471564
rect 580073 471472 584960 471474
rect 580073 471416 580078 471472
rect 580134 471416 584960 471472
rect 580073 471414 584960 471416
rect 580073 471411 580139 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580901 458146 580967 458149
rect 583520 458146 584960 458236
rect 580901 458144 584960 458146
rect 580901 458088 580906 458144
rect 580962 458088 584960 458144
rect 580901 458086 584960 458088
rect 580901 458083 580967 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580809 431626 580875 431629
rect 583520 431626 584960 431716
rect 580809 431624 584960 431626
rect 580809 431568 580814 431624
rect 580870 431568 584960 431624
rect 580809 431566 584960 431568
rect 580809 431563 580875 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3693 397490 3759 397493
rect -960 397488 3759 397490
rect -960 397432 3698 397488
rect 3754 397432 3759 397488
rect -960 397430 3759 397432
rect -960 397340 480 397430
rect 3693 397427 3759 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 4061 358458 4127 358461
rect -960 358456 4127 358458
rect -960 358400 4066 358456
rect 4122 358400 4127 358456
rect -960 358398 4127 358400
rect -960 358308 480 358398
rect 4061 358395 4127 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3877 345402 3943 345405
rect -960 345400 3943 345402
rect -960 345344 3882 345400
rect 3938 345344 3943 345400
rect -960 345342 3943 345344
rect -960 345252 480 345342
rect 3877 345339 3943 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579981 298754 580047 298757
rect 583520 298754 584960 298844
rect 579981 298752 584960 298754
rect 579981 298696 579986 298752
rect 580042 298696 584960 298752
rect 579981 298694 584960 298696
rect 579981 298691 580047 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579981 272234 580047 272237
rect 583520 272234 584960 272324
rect 579981 272232 584960 272234
rect 579981 272176 579986 272232
rect 580042 272176 584960 272232
rect 579981 272174 584960 272176
rect 579981 272171 580047 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3141 267202 3207 267205
rect -960 267200 3207 267202
rect -960 267144 3146 267200
rect 3202 267144 3207 267200
rect -960 267142 3207 267144
rect -960 267052 480 267142
rect 3141 267139 3207 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3233 254146 3299 254149
rect -960 254144 3299 254146
rect -960 254088 3238 254144
rect 3294 254088 3299 254144
rect -960 254086 3299 254088
rect -960 253996 480 254086
rect 3233 254083 3299 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3233 228034 3299 228037
rect -960 228032 3299 228034
rect -960 227976 3238 228032
rect 3294 227976 3299 228032
rect -960 227974 3299 227976
rect -960 227884 480 227974
rect 3233 227971 3299 227974
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3233 214978 3299 214981
rect -960 214976 3299 214978
rect -960 214920 3238 214976
rect 3294 214920 3299 214976
rect -960 214918 3299 214920
rect -960 214828 480 214918
rect 3233 214915 3299 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 140773 195666 140839 195669
rect 143582 195666 144164 195674
rect 140773 195664 144164 195666
rect 140773 195608 140778 195664
rect 140834 195614 144164 195664
rect 140834 195608 143642 195614
rect 140773 195606 143642 195608
rect 140773 195603 140839 195606
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 149605 193354 149671 193357
rect 165429 193354 165495 193357
rect 149605 193352 165495 193354
rect 149605 193296 149610 193352
rect 149666 193296 165434 193352
rect 165490 193296 165495 193352
rect 149605 193294 165495 193296
rect 149605 193291 149671 193294
rect 165429 193291 165495 193294
rect 579797 192538 579863 192541
rect 583520 192538 584960 192628
rect 579797 192536 584960 192538
rect 579797 192480 579802 192536
rect 579858 192480 584960 192536
rect 579797 192478 584960 192480
rect 579797 192475 579863 192478
rect 583520 192388 584960 192478
rect 140773 191858 140839 191861
rect 143214 191858 143980 191900
rect 140773 191856 143980 191858
rect 140773 191800 140778 191856
rect 140834 191840 143980 191856
rect 140834 191800 143274 191840
rect 140773 191798 143274 191800
rect 140773 191795 140839 191798
rect 140957 191722 141023 191725
rect 143398 191722 143980 191760
rect 140957 191720 143980 191722
rect 140957 191664 140962 191720
rect 141018 191700 143980 191720
rect 141018 191664 143458 191700
rect 140957 191662 143458 191664
rect 140957 191659 141023 191662
rect 140865 191586 140931 191589
rect 143582 191586 144164 191630
rect 140865 191584 144164 191586
rect 140865 191528 140870 191584
rect 140926 191570 144164 191584
rect 140926 191528 143642 191570
rect 140865 191526 143642 191528
rect 140865 191523 140931 191526
rect 140773 190906 140839 190909
rect 144134 190906 144194 191460
rect 140773 190904 144194 190906
rect 140773 190848 140778 190904
rect 140834 190848 144194 190904
rect 140773 190846 144194 190848
rect 140773 190843 140839 190846
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 139393 187642 139459 187645
rect 144126 187642 144132 187644
rect 139393 187640 144132 187642
rect 139393 187584 139398 187640
rect 139454 187584 144132 187640
rect 139393 187582 144132 187584
rect 139393 187579 139459 187582
rect 144126 187580 144132 187582
rect 144196 187580 144202 187644
rect 140773 186284 140839 186285
rect 140773 186282 140820 186284
rect 140728 186280 140820 186282
rect 140728 186224 140778 186280
rect 140728 186222 140820 186224
rect 140773 186220 140820 186222
rect 140884 186220 140890 186284
rect 140773 186219 140839 186220
rect 140957 182746 141023 182749
rect 143022 182746 143028 182748
rect 140957 182744 143028 182746
rect 140957 182688 140962 182744
rect 141018 182688 143028 182744
rect 140957 182686 143028 182688
rect 140957 182683 141023 182686
rect 143022 182684 143028 182686
rect 143092 182684 143098 182748
rect 140773 182610 140839 182613
rect 141550 182610 141556 182612
rect 140773 182608 141556 182610
rect 140773 182552 140778 182608
rect 140834 182552 141556 182608
rect 140773 182550 141556 182552
rect 140773 182547 140839 182550
rect 141550 182548 141556 182550
rect 141620 182548 141626 182612
rect 140865 182474 140931 182477
rect 140998 182474 141004 182476
rect 140865 182472 141004 182474
rect 140865 182416 140870 182472
rect 140926 182416 141004 182472
rect 140865 182414 141004 182416
rect 140865 182411 140931 182414
rect 140998 182412 141004 182414
rect 141068 182412 141074 182476
rect 142470 180916 142476 180980
rect 142540 180978 142546 180980
rect 144637 180978 144703 180981
rect 142540 180976 144703 180978
rect 142540 180920 144642 180976
rect 144698 180920 144703 180976
rect 142540 180918 144703 180920
rect 142540 180916 142546 180918
rect 144637 180915 144703 180918
rect 146017 180978 146083 180981
rect 146150 180978 146156 180980
rect 146017 180976 146156 180978
rect 146017 180920 146022 180976
rect 146078 180920 146156 180976
rect 146017 180918 146156 180920
rect 146017 180915 146083 180918
rect 146150 180916 146156 180918
rect 146220 180916 146226 180980
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect 143022 178876 143028 178940
rect 143092 178938 143098 178940
rect 144085 178938 144151 178941
rect 143092 178936 144151 178938
rect 143092 178880 144090 178936
rect 144146 178880 144151 178936
rect 143092 178878 144151 178880
rect 143092 178876 143098 178878
rect 144085 178875 144151 178878
rect 140998 178740 141004 178804
rect 141068 178802 141074 178804
rect 141601 178802 141667 178805
rect 141068 178800 141667 178802
rect 141068 178744 141606 178800
rect 141662 178744 141667 178800
rect 141068 178742 141667 178744
rect 141068 178740 141074 178742
rect 141601 178739 141667 178742
rect 140814 178604 140820 178668
rect 140884 178666 140890 178668
rect 142061 178666 142127 178669
rect 140884 178664 142127 178666
rect 140884 178608 142066 178664
rect 142122 178608 142127 178664
rect 140884 178606 142127 178608
rect 140884 178604 140890 178606
rect 142061 178603 142127 178606
rect 141550 178468 141556 178532
rect 141620 178530 141626 178532
rect 141693 178530 141759 178533
rect 141620 178528 141759 178530
rect 141620 178472 141698 178528
rect 141754 178472 141759 178528
rect 141620 178470 141759 178472
rect 141620 178468 141626 178470
rect 141693 178467 141759 178470
rect -960 175796 480 176036
rect 165429 175540 165495 175541
rect 165429 175536 165476 175540
rect 165540 175538 165546 175540
rect 165429 175480 165434 175536
rect 165429 175476 165476 175480
rect 165540 175478 165586 175538
rect 165540 175476 165546 175478
rect 165429 175475 165495 175476
rect 149329 175402 149395 175405
rect 154389 175402 154455 175405
rect 149329 175400 154455 175402
rect 149329 175344 149334 175400
rect 149390 175344 154394 175400
rect 154450 175344 154455 175400
rect 149329 175342 154455 175344
rect 149329 175339 149395 175342
rect 154389 175339 154455 175342
rect 146150 174524 146156 174588
rect 146220 174586 146226 174588
rect 171133 174586 171199 174589
rect 146220 174584 171199 174586
rect 146220 174528 171138 174584
rect 171194 174528 171199 174584
rect 146220 174526 171199 174528
rect 146220 174524 146226 174526
rect 171133 174523 171199 174526
rect 142521 172956 142587 172957
rect 142470 172954 142476 172956
rect 142430 172894 142476 172954
rect 142540 172952 142587 172956
rect 165429 172956 165495 172957
rect 165429 172954 165476 172956
rect 142582 172896 142587 172952
rect 142470 172892 142476 172894
rect 142540 172892 142587 172896
rect 165384 172952 165476 172954
rect 165384 172896 165434 172952
rect 165384 172894 165476 172896
rect 142521 172891 142587 172892
rect 165429 172892 165476 172894
rect 165540 172892 165546 172956
rect 165429 172891 165495 172892
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3141 162890 3207 162893
rect -960 162888 3207 162890
rect -960 162832 3146 162888
rect 3202 162832 3207 162888
rect -960 162830 3207 162832
rect -960 162740 480 162830
rect 3141 162827 3207 162830
rect 144126 156572 144132 156636
rect 144196 156634 144202 156636
rect 155217 156634 155283 156637
rect 144196 156632 155283 156634
rect 144196 156576 155222 156632
rect 155278 156576 155283 156632
rect 144196 156574 155283 156576
rect 144196 156572 144202 156574
rect 155217 156571 155283 156574
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 45001 141402 45067 141405
rect 182214 141402 182220 141404
rect 45001 141400 182220 141402
rect 45001 141344 45006 141400
rect 45062 141344 182220 141400
rect 45001 141342 182220 141344
rect 45001 141339 45067 141342
rect 182214 141340 182220 141342
rect 182284 141340 182290 141404
rect 118550 139980 118556 140044
rect 118620 140042 118626 140044
rect 580441 140042 580507 140045
rect 118620 140040 580507 140042
rect 118620 139984 580446 140040
rect 580502 139984 580507 140040
rect 118620 139982 580507 139984
rect 118620 139980 118626 139982
rect 580441 139979 580507 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 118417 136642 118483 136645
rect 118417 136640 120060 136642
rect 118417 136584 118422 136640
rect 118478 136584 120060 136640
rect 118417 136582 120060 136584
rect 118417 136579 118483 136582
rect 118233 136098 118299 136101
rect 120625 136098 120691 136101
rect 118233 136096 120691 136098
rect 118233 136040 118238 136096
rect 118294 136040 120630 136096
rect 120686 136040 120691 136096
rect 118233 136038 120691 136040
rect 118233 136035 118299 136038
rect 120582 136035 120691 136038
rect 120582 135524 120642 136035
rect 118417 135010 118483 135013
rect 120533 135010 120599 135013
rect 118417 135008 120642 135010
rect 118417 134952 118422 135008
rect 118478 134952 120538 135008
rect 120594 134952 120642 135008
rect 118417 134950 120642 134952
rect 118417 134947 118483 134950
rect 120533 134947 120642 134950
rect 120582 134436 120642 134947
rect 117313 133378 117379 133381
rect 117313 133376 120060 133378
rect 117313 133320 117318 133376
rect 117374 133320 120060 133376
rect 117313 133318 120060 133320
rect 117313 133315 117379 133318
rect 116945 132290 117011 132293
rect 116945 132288 120060 132290
rect 116945 132232 116950 132288
rect 117006 132232 120060 132288
rect 116945 132230 120060 132232
rect 116945 132227 117011 132230
rect 116853 131202 116919 131205
rect 116853 131200 120060 131202
rect 116853 131144 116858 131200
rect 116914 131144 120060 131200
rect 116853 131142 120060 131144
rect 116853 131139 116919 131142
rect 181069 131066 181135 131069
rect 179860 131064 181135 131066
rect 179860 131008 181074 131064
rect 181130 131008 181135 131064
rect 179860 131006 181135 131008
rect 181069 131003 181135 131006
rect 116669 130114 116735 130117
rect 116669 130112 120060 130114
rect 116669 130056 116674 130112
rect 116730 130056 120060 130112
rect 116669 130054 120060 130056
rect 116669 130051 116735 130054
rect 180885 129706 180951 129709
rect 179860 129704 180951 129706
rect 179860 129648 180890 129704
rect 180946 129648 180951 129704
rect 179860 129646 180951 129648
rect 180885 129643 180951 129646
rect 117313 129026 117379 129029
rect 117313 129024 120060 129026
rect 117313 128968 117318 129024
rect 117374 128968 120060 129024
rect 117313 128966 120060 128968
rect 117313 128963 117379 128966
rect 179462 128213 179522 128316
rect 179462 128208 179571 128213
rect 179462 128152 179510 128208
rect 179566 128152 179571 128208
rect 179462 128150 179571 128152
rect 179505 128147 179571 128150
rect 117313 127938 117379 127941
rect 117313 127936 120060 127938
rect 117313 127880 117318 127936
rect 117374 127880 120060 127936
rect 117313 127878 120060 127880
rect 117313 127875 117379 127878
rect 179462 126853 179522 126956
rect 117681 126850 117747 126853
rect 117681 126848 120060 126850
rect 117681 126792 117686 126848
rect 117742 126792 120060 126848
rect 117681 126790 120060 126792
rect 179413 126848 179522 126853
rect 179413 126792 179418 126848
rect 179474 126792 179522 126848
rect 179413 126790 179522 126792
rect 117681 126787 117747 126790
rect 179413 126787 179479 126790
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 117313 125762 117379 125765
rect 117865 125762 117931 125765
rect 117313 125760 120060 125762
rect 117313 125704 117318 125760
rect 117374 125704 117870 125760
rect 117926 125704 120060 125760
rect 117313 125702 120060 125704
rect 117313 125699 117379 125702
rect 117865 125699 117931 125702
rect 180793 125626 180859 125629
rect 179860 125624 180859 125626
rect 179860 125568 180798 125624
rect 180854 125568 180859 125624
rect 179860 125566 180859 125568
rect 180793 125563 180859 125566
rect -960 123572 480 123812
rect 117773 123586 117839 123589
rect 120030 123586 120090 124644
rect 182173 124266 182239 124269
rect 179860 124264 182239 124266
rect 179860 124208 182178 124264
rect 182234 124208 182239 124264
rect 179860 124206 182239 124208
rect 182173 124203 182239 124206
rect 117773 123584 120090 123586
rect 117773 123528 117778 123584
rect 117834 123556 120090 123584
rect 117834 123528 120060 123556
rect 117773 123526 120060 123528
rect 117773 123523 117839 123526
rect 183001 122906 183067 122909
rect 179860 122904 183067 122906
rect 179860 122848 183006 122904
rect 183062 122848 183067 122904
rect 179860 122846 183067 122848
rect 183001 122843 183067 122846
rect 117681 122498 117747 122501
rect 117681 122496 120060 122498
rect 117681 122440 117686 122496
rect 117742 122440 120060 122496
rect 117681 122438 120060 122440
rect 117681 122435 117747 122438
rect 182909 121546 182975 121549
rect 179860 121544 182975 121546
rect 179860 121488 182914 121544
rect 182970 121488 182975 121544
rect 179860 121486 182975 121488
rect 182909 121483 182975 121486
rect 117405 121410 117471 121413
rect 117405 121408 120060 121410
rect 117405 121352 117410 121408
rect 117466 121352 120060 121408
rect 117405 121350 120060 121352
rect 117405 121347 117471 121350
rect 117313 120322 117379 120325
rect 117313 120320 120060 120322
rect 117313 120264 117318 120320
rect 117374 120264 120060 120320
rect 117313 120262 120060 120264
rect 117313 120259 117379 120262
rect 182725 120186 182791 120189
rect 179860 120184 182791 120186
rect 179860 120128 182730 120184
rect 182786 120128 182791 120184
rect 179860 120126 182791 120128
rect 182725 120123 182791 120126
rect 117865 119234 117931 119237
rect 117865 119232 120060 119234
rect 117865 119176 117870 119232
rect 117926 119176 120060 119232
rect 117865 119174 120060 119176
rect 117865 119171 117931 119174
rect 182633 118826 182699 118829
rect 179860 118824 182699 118826
rect 179860 118768 182638 118824
rect 182694 118768 182699 118824
rect 179860 118766 182699 118768
rect 182633 118763 182699 118766
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 182541 117466 182607 117469
rect 179860 117464 182607 117466
rect 179860 117408 182546 117464
rect 182602 117408 182607 117464
rect 179860 117406 182607 117408
rect 182541 117403 182607 117406
rect 117313 117058 117379 117061
rect 117313 117056 120060 117058
rect 117313 117000 117318 117056
rect 117374 117000 120060 117056
rect 117313 116998 120060 117000
rect 117313 116995 117379 116998
rect 182449 116106 182515 116109
rect 179860 116104 182515 116106
rect 179860 116048 182454 116104
rect 182510 116048 182515 116104
rect 179860 116046 182515 116048
rect 182449 116043 182515 116046
rect 117405 115970 117471 115973
rect 117405 115968 120060 115970
rect 117405 115912 117410 115968
rect 117466 115912 120060 115968
rect 117405 115910 120060 115912
rect 117405 115907 117471 115910
rect 117313 114882 117379 114885
rect 117313 114880 120060 114882
rect 117313 114824 117318 114880
rect 117374 114824 120060 114880
rect 117313 114822 120060 114824
rect 117313 114819 117379 114822
rect 182357 114746 182423 114749
rect 179860 114744 182423 114746
rect 179860 114688 182362 114744
rect 182418 114688 182423 114744
rect 179860 114686 182423 114688
rect 182357 114683 182423 114686
rect 117313 113794 117379 113797
rect 117313 113792 120060 113794
rect 117313 113736 117318 113792
rect 117374 113736 120060 113792
rect 117313 113734 120060 113736
rect 117313 113731 117379 113734
rect 182265 113386 182331 113389
rect 179860 113384 182331 113386
rect 179860 113328 182270 113384
rect 182326 113328 182331 113384
rect 179860 113326 182331 113328
rect 182265 113323 182331 113326
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 117313 112706 117379 112709
rect 117313 112704 120060 112706
rect 117313 112648 117318 112704
rect 117374 112648 120060 112704
rect 583520 112692 584960 112782
rect 117313 112646 120060 112648
rect 117313 112643 117379 112646
rect 182817 112026 182883 112029
rect 179860 112024 182883 112026
rect 179860 111968 182822 112024
rect 182878 111968 182883 112024
rect 179860 111966 182883 111968
rect 182817 111963 182883 111966
rect 117313 111618 117379 111621
rect 117313 111616 120060 111618
rect 117313 111560 117318 111616
rect 117374 111560 120060 111616
rect 117313 111558 120060 111560
rect 117313 111555 117379 111558
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect 182214 110666 182220 110668
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect 179860 110606 182220 110666
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 182214 110604 182220 110606
rect 182284 110604 182290 110668
rect 117405 110530 117471 110533
rect 117405 110528 120060 110530
rect 117405 110472 117410 110528
rect 117466 110472 120060 110528
rect 117405 110470 120060 110472
rect 117405 110467 117471 110470
rect 117313 109442 117379 109445
rect 117313 109440 120060 109442
rect 117313 109384 117318 109440
rect 117374 109384 120060 109440
rect 117313 109382 120060 109384
rect 117313 109379 117379 109382
rect 182173 109306 182239 109309
rect 179860 109304 182239 109306
rect 179860 109248 182178 109304
rect 182234 109248 182239 109304
rect 179860 109246 182239 109248
rect 182173 109243 182239 109246
rect 117313 108354 117379 108357
rect 117313 108352 120060 108354
rect 117313 108296 117318 108352
rect 117374 108296 120060 108352
rect 117313 108294 120060 108296
rect 117313 108291 117379 108294
rect 180977 107946 181043 107949
rect 179860 107944 181043 107946
rect 179860 107888 180982 107944
rect 181038 107888 181043 107944
rect 179860 107886 181043 107888
rect 180977 107883 181043 107886
rect 117313 107266 117379 107269
rect 117313 107264 120060 107266
rect 117313 107208 117318 107264
rect 117374 107208 120060 107264
rect 117313 107206 120060 107208
rect 117313 107203 117379 107206
rect 183277 106586 183343 106589
rect 179860 106584 183343 106586
rect 179860 106528 183282 106584
rect 183338 106528 183343 106584
rect 179860 106526 183343 106528
rect 183277 106523 183343 106526
rect 117313 106178 117379 106181
rect 117313 106176 120060 106178
rect 117313 106120 117318 106176
rect 117374 106120 120060 106176
rect 117313 106118 120060 106120
rect 117313 106115 117379 106118
rect 183277 105226 183343 105229
rect 179860 105224 183343 105226
rect 179860 105168 183282 105224
rect 183338 105168 183343 105224
rect 179860 105166 183343 105168
rect 183277 105163 183343 105166
rect 117405 105090 117471 105093
rect 117405 105088 120060 105090
rect 117405 105032 117410 105088
rect 117466 105032 120060 105088
rect 117405 105030 120060 105032
rect 117405 105027 117471 105030
rect 117313 104002 117379 104005
rect 117313 104000 120060 104002
rect 117313 103944 117318 104000
rect 117374 103944 120060 104000
rect 117313 103942 120060 103944
rect 117313 103939 117379 103942
rect 183277 103866 183343 103869
rect 179860 103864 183343 103866
rect 179860 103808 183282 103864
rect 183338 103808 183343 103864
rect 179860 103806 183343 103808
rect 183277 103803 183343 103806
rect 118601 102914 118667 102917
rect 118601 102912 120060 102914
rect 118601 102856 118606 102912
rect 118662 102856 120060 102912
rect 118601 102854 120060 102856
rect 118601 102851 118667 102854
rect 183277 102506 183343 102509
rect 179860 102504 183343 102506
rect 179860 102448 183282 102504
rect 183338 102448 183343 102504
rect 179860 102446 183343 102448
rect 183277 102443 183343 102446
rect 119153 101826 119219 101829
rect 119153 101824 120060 101826
rect 119153 101768 119158 101824
rect 119214 101768 120060 101824
rect 119153 101766 120060 101768
rect 119153 101763 119219 101766
rect 183277 101146 183343 101149
rect 179860 101144 183343 101146
rect 179860 101088 183282 101144
rect 183338 101088 183343 101144
rect 179860 101086 183343 101088
rect 183277 101083 183343 101086
rect 119245 100738 119311 100741
rect 119245 100736 120060 100738
rect 119245 100680 119250 100736
rect 119306 100680 120060 100736
rect 119245 100678 120060 100680
rect 119245 100675 119311 100678
rect 183185 99786 183251 99789
rect 179860 99784 183251 99786
rect 179860 99728 183190 99784
rect 183246 99728 183251 99784
rect 179860 99726 183251 99728
rect 183185 99723 183251 99726
rect 119061 99650 119127 99653
rect 119061 99648 120060 99650
rect 119061 99592 119066 99648
rect 119122 99592 120060 99648
rect 119061 99590 120060 99592
rect 119061 99587 119127 99590
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 118969 98562 119035 98565
rect 118969 98560 120060 98562
rect 118969 98504 118974 98560
rect 119030 98504 120060 98560
rect 118969 98502 120060 98504
rect 118969 98499 119035 98502
rect 183185 98426 183251 98429
rect 179860 98424 183251 98426
rect 179860 98368 183190 98424
rect 183246 98368 183251 98424
rect 179860 98366 183251 98368
rect 183185 98363 183251 98366
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 118877 97474 118943 97477
rect 118877 97472 120060 97474
rect 118877 97416 118882 97472
rect 118938 97416 120060 97472
rect 118877 97414 120060 97416
rect 118877 97411 118943 97414
rect 183185 97066 183251 97069
rect 179860 97064 183251 97066
rect 179860 97008 183190 97064
rect 183246 97008 183251 97064
rect 179860 97006 183251 97008
rect 183185 97003 183251 97006
rect 118550 96324 118556 96388
rect 118620 96386 118626 96388
rect 118620 96326 120060 96386
rect 118620 96324 118626 96326
rect 183185 95706 183251 95709
rect 179860 95704 183251 95706
rect 179860 95648 183190 95704
rect 183246 95648 183251 95704
rect 179860 95646 183251 95648
rect 183185 95643 183251 95646
rect 118785 95298 118851 95301
rect 118785 95296 120060 95298
rect 118785 95240 118790 95296
rect 118846 95240 120060 95296
rect 118785 95238 120060 95240
rect 118785 95235 118851 95238
rect 183461 94346 183527 94349
rect 179860 94344 183527 94346
rect 179860 94288 183466 94344
rect 183522 94288 183527 94344
rect 179860 94286 183527 94288
rect 183461 94283 183527 94286
rect 118049 94210 118115 94213
rect 118049 94208 120060 94210
rect 118049 94152 118054 94208
rect 118110 94152 120060 94208
rect 118049 94150 120060 94152
rect 118049 94147 118115 94150
rect 118325 93122 118391 93125
rect 118325 93120 120060 93122
rect 118325 93064 118330 93120
rect 118386 93064 120060 93120
rect 118325 93062 120060 93064
rect 118325 93059 118391 93062
rect 183461 92986 183527 92989
rect 179860 92984 183527 92986
rect 179860 92928 183466 92984
rect 183522 92928 183527 92984
rect 179860 92926 183527 92928
rect 183461 92923 183527 92926
rect 118141 92034 118207 92037
rect 118141 92032 120060 92034
rect 118141 91976 118146 92032
rect 118202 91976 120060 92032
rect 118141 91974 120060 91976
rect 118141 91971 118207 91974
rect 183461 91626 183527 91629
rect 179860 91624 183527 91626
rect 179860 91568 183466 91624
rect 183522 91568 183527 91624
rect 179860 91566 183527 91568
rect 183461 91563 183527 91566
rect 118233 90946 118299 90949
rect 118233 90944 120060 90946
rect 118233 90888 118238 90944
rect 118294 90888 120060 90944
rect 118233 90886 120060 90888
rect 118233 90883 118299 90886
rect 183461 90266 183527 90269
rect 179860 90264 183527 90266
rect 179860 90208 183466 90264
rect 183522 90208 183527 90264
rect 179860 90206 183527 90208
rect 183461 90203 183527 90206
rect 118417 89858 118483 89861
rect 118417 89856 120060 89858
rect 118417 89800 118422 89856
rect 118478 89800 120060 89856
rect 118417 89798 120060 89800
rect 118417 89795 118483 89798
rect 182265 88906 182331 88909
rect 179860 88904 182331 88906
rect 179860 88848 182270 88904
rect 182326 88848 182331 88904
rect 179860 88846 182331 88848
rect 182265 88843 182331 88846
rect 118693 88770 118759 88773
rect 118693 88768 120060 88770
rect 118693 88712 118698 88768
rect 118754 88712 120060 88768
rect 118693 88710 120060 88712
rect 118693 88707 118759 88710
rect 118509 87682 118575 87685
rect 118509 87680 120060 87682
rect 118509 87624 118514 87680
rect 118570 87624 120060 87680
rect 118509 87622 120060 87624
rect 118509 87619 118575 87622
rect 182817 87546 182883 87549
rect 179860 87544 182883 87546
rect 179860 87488 182822 87544
rect 182878 87488 182883 87544
rect 179860 87486 182883 87488
rect 182817 87483 182883 87486
rect 118509 86594 118575 86597
rect 118509 86592 120060 86594
rect 118509 86536 118514 86592
rect 118570 86536 120060 86592
rect 118509 86534 120060 86536
rect 118509 86531 118575 86534
rect 182725 86186 182791 86189
rect 179860 86184 182791 86186
rect 179860 86128 182730 86184
rect 182786 86128 182791 86184
rect 179860 86126 182791 86128
rect 182725 86123 182791 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 118601 85506 118667 85509
rect 118601 85504 120060 85506
rect 118601 85448 118606 85504
rect 118662 85448 120060 85504
rect 118601 85446 120060 85448
rect 118601 85443 118667 85446
rect 182725 84826 182791 84829
rect 179860 84824 182791 84826
rect -960 84690 480 84780
rect 179860 84768 182730 84824
rect 182786 84768 182791 84824
rect 179860 84766 182791 84768
rect 182725 84763 182791 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 118233 84418 118299 84421
rect 118233 84416 120060 84418
rect 118233 84360 118238 84416
rect 118294 84360 120060 84416
rect 118233 84358 120060 84360
rect 118233 84355 118299 84358
rect 182725 83466 182791 83469
rect 179860 83464 182791 83466
rect 179860 83408 182730 83464
rect 182786 83408 182791 83464
rect 179860 83406 182791 83408
rect 182725 83403 182791 83406
rect 118325 83330 118391 83333
rect 118325 83328 120060 83330
rect 118325 83272 118330 83328
rect 118386 83272 120060 83328
rect 118325 83270 120060 83272
rect 118325 83267 118391 83270
rect 182909 82106 182975 82109
rect 179860 82104 182975 82106
rect 179860 82048 182914 82104
rect 182970 82048 182975 82104
rect 179860 82046 182975 82048
rect 182909 82043 182975 82046
rect 182817 80746 182883 80749
rect 179860 80744 182883 80746
rect 179860 80688 182822 80744
rect 182878 80688 182883 80744
rect 179860 80686 182883 80688
rect 182817 80683 182883 80686
rect 171358 80548 171364 80612
rect 171428 80610 171434 80612
rect 393957 80610 394023 80613
rect 171428 80608 394023 80610
rect 171428 80552 393962 80608
rect 394018 80552 394023 80608
rect 171428 80550 394023 80552
rect 171428 80548 171434 80550
rect 393957 80547 394023 80550
rect 44909 80474 44975 80477
rect 44909 80472 173220 80474
rect 44909 80416 44914 80472
rect 44970 80416 173220 80472
rect 44909 80414 173220 80416
rect 44909 80411 44975 80414
rect 172278 80338 172284 80340
rect 164558 80278 172284 80338
rect 125225 80202 125291 80205
rect 125225 80200 133016 80202
rect 125225 80144 125230 80200
rect 125286 80144 133016 80200
rect 125225 80142 133016 80144
rect 125225 80139 125291 80142
rect 129774 80066 129780 80068
rect 129736 80004 129780 80066
rect 129844 80004 129850 80068
rect 126743 79964 126809 79967
rect 126700 79962 126809 79964
rect 124765 79930 124831 79933
rect 126099 79930 126165 79933
rect 124765 79928 126165 79930
rect 124765 79872 124770 79928
rect 124826 79872 126104 79928
rect 126160 79872 126165 79928
rect 124765 79870 126165 79872
rect 124765 79867 124831 79870
rect 126099 79867 126165 79870
rect 126278 79868 126284 79932
rect 126348 79930 126354 79932
rect 126559 79930 126625 79933
rect 126348 79928 126625 79930
rect 126348 79872 126564 79928
rect 126620 79872 126625 79928
rect 126348 79870 126625 79872
rect 126348 79868 126354 79870
rect 126559 79867 126625 79870
rect 126700 79906 126748 79962
rect 126804 79906 126809 79962
rect 126700 79901 126809 79906
rect 127111 79962 127177 79967
rect 127111 79906 127116 79962
rect 127172 79906 127177 79962
rect 127111 79901 127177 79906
rect 127295 79964 127361 79967
rect 127295 79962 127404 79964
rect 127295 79906 127300 79962
rect 127356 79932 127404 79962
rect 127755 79962 127821 79967
rect 127356 79906 127388 79932
rect 127295 79901 127388 79906
rect 125317 79794 125383 79797
rect 126700 79794 126760 79901
rect 125317 79792 126760 79794
rect 125317 79736 125322 79792
rect 125378 79736 126760 79792
rect 125317 79734 126760 79736
rect 127114 79794 127174 79901
rect 127344 79870 127388 79901
rect 127382 79868 127388 79870
rect 127452 79868 127458 79932
rect 127571 79928 127637 79933
rect 127755 79932 127760 79962
rect 127816 79932 127821 79962
rect 127571 79872 127576 79928
rect 127632 79872 127637 79928
rect 127571 79867 127637 79872
rect 127750 79868 127756 79932
rect 127820 79930 127826 79932
rect 128307 79930 128373 79933
rect 127820 79870 127878 79930
rect 128126 79928 128373 79930
rect 128126 79872 128312 79928
rect 128368 79872 128373 79928
rect 128126 79870 128373 79872
rect 127820 79868 127826 79870
rect 127382 79794 127388 79796
rect 127114 79734 127388 79794
rect 125317 79731 125383 79734
rect 127382 79732 127388 79734
rect 127452 79732 127458 79796
rect 127574 79658 127634 79867
rect 127985 79658 128051 79661
rect 127574 79656 128051 79658
rect 127574 79600 127990 79656
rect 128046 79600 128051 79656
rect 127574 79598 128051 79600
rect 128126 79658 128186 79870
rect 128307 79867 128373 79870
rect 128486 79868 128492 79932
rect 128556 79930 128562 79932
rect 128675 79930 128741 79933
rect 129227 79932 129293 79933
rect 128556 79928 128741 79930
rect 128556 79872 128680 79928
rect 128736 79872 128741 79928
rect 128556 79870 128741 79872
rect 128556 79868 128562 79870
rect 128675 79867 128741 79870
rect 129222 79868 129228 79932
rect 129292 79930 129298 79932
rect 129736 79930 129796 80004
rect 132956 79967 133016 80142
rect 140998 80140 141004 80204
rect 141068 80202 141074 80204
rect 144862 80202 144868 80204
rect 141068 80142 142170 80202
rect 141068 80140 141074 80142
rect 142110 79967 142170 80142
rect 142938 80142 144868 80202
rect 142938 79967 142998 80142
rect 144862 80140 144868 80142
rect 144932 80140 144938 80204
rect 152406 80140 152412 80204
rect 152476 80202 152482 80204
rect 152476 80142 152934 80202
rect 152476 80140 152482 80142
rect 145414 80066 145420 80068
rect 144870 80006 145420 80066
rect 131159 79962 131225 79967
rect 129871 79930 129937 79933
rect 129292 79870 129384 79930
rect 129736 79928 129937 79930
rect 129736 79872 129876 79928
rect 129932 79872 129937 79928
rect 129736 79870 129937 79872
rect 129292 79868 129298 79870
rect 129227 79867 129293 79868
rect 129871 79867 129937 79870
rect 130055 79930 130121 79933
rect 130055 79928 130394 79930
rect 130055 79872 130060 79928
rect 130116 79872 130394 79928
rect 130055 79870 130394 79872
rect 130055 79867 130121 79870
rect 130334 79796 130394 79870
rect 130878 79868 130884 79932
rect 130948 79930 130954 79932
rect 131159 79930 131164 79962
rect 130948 79906 131164 79930
rect 131220 79906 131225 79962
rect 132171 79962 132237 79967
rect 130948 79901 131225 79906
rect 131343 79930 131409 79933
rect 132171 79932 132176 79962
rect 132232 79932 132237 79962
rect 132539 79962 132605 79967
rect 131343 79928 131682 79930
rect 130948 79870 131222 79901
rect 131343 79872 131348 79928
rect 131404 79872 131682 79928
rect 131343 79870 131682 79872
rect 130948 79868 130954 79870
rect 131343 79867 131409 79870
rect 130326 79732 130332 79796
rect 130396 79732 130402 79796
rect 128261 79658 128327 79661
rect 128721 79660 128787 79661
rect 128670 79658 128676 79660
rect 128126 79656 128327 79658
rect 128126 79600 128266 79656
rect 128322 79600 128327 79656
rect 128126 79598 128327 79600
rect 128630 79598 128676 79658
rect 128740 79656 128787 79660
rect 128782 79600 128787 79656
rect 127985 79595 128051 79598
rect 128261 79595 128327 79598
rect 128670 79596 128676 79598
rect 128740 79596 128787 79600
rect 131246 79596 131252 79660
rect 131316 79658 131322 79660
rect 131622 79658 131682 79870
rect 132166 79868 132172 79932
rect 132236 79930 132242 79932
rect 132236 79870 132294 79930
rect 132539 79906 132544 79962
rect 132600 79906 132605 79962
rect 132539 79901 132605 79906
rect 132956 79962 133065 79967
rect 134471 79964 134537 79967
rect 132956 79906 133004 79962
rect 133060 79906 133065 79962
rect 134428 79962 134537 79964
rect 132956 79904 133065 79906
rect 132999 79901 133065 79904
rect 132236 79868 132242 79870
rect 132542 79794 132602 79901
rect 133454 79868 133460 79932
rect 133524 79930 133530 79932
rect 133919 79930 133985 79933
rect 134287 79930 134353 79933
rect 133524 79928 133985 79930
rect 133524 79872 133924 79928
rect 133980 79872 133985 79928
rect 133524 79870 133985 79872
rect 133524 79868 133530 79870
rect 133919 79867 133985 79870
rect 134152 79928 134353 79930
rect 134152 79872 134292 79928
rect 134348 79872 134353 79928
rect 134152 79870 134353 79872
rect 132769 79794 132835 79797
rect 132542 79792 132835 79794
rect 132542 79736 132774 79792
rect 132830 79736 132835 79792
rect 132542 79734 132835 79736
rect 132769 79731 132835 79734
rect 131316 79598 131682 79658
rect 132677 79658 132743 79661
rect 133086 79658 133092 79660
rect 132677 79656 133092 79658
rect 132677 79600 132682 79656
rect 132738 79600 133092 79656
rect 132677 79598 133092 79600
rect 131316 79596 131322 79598
rect 128721 79595 128787 79596
rect 132677 79595 132743 79598
rect 133086 79596 133092 79598
rect 133156 79596 133162 79660
rect 134152 79658 134212 79870
rect 134287 79867 134353 79870
rect 134428 79906 134476 79962
rect 134532 79906 134537 79962
rect 134931 79962 134997 79967
rect 136495 79964 136561 79967
rect 134428 79901 134537 79906
rect 134747 79928 134813 79933
rect 134428 79797 134488 79901
rect 134747 79872 134752 79928
rect 134808 79872 134813 79928
rect 134931 79906 134936 79962
rect 134992 79906 134997 79962
rect 136222 79962 136561 79964
rect 134931 79901 134997 79906
rect 135391 79930 135457 79933
rect 135391 79928 135500 79930
rect 134747 79867 134813 79872
rect 134425 79792 134491 79797
rect 134425 79736 134430 79792
rect 134486 79736 134491 79792
rect 134425 79731 134491 79736
rect 134750 79661 134810 79867
rect 134934 79797 134994 79901
rect 135391 79872 135396 79928
rect 135452 79872 135500 79928
rect 135391 79867 135500 79872
rect 135667 79928 135733 79933
rect 135667 79872 135672 79928
rect 135728 79872 135733 79928
rect 135667 79867 135733 79872
rect 136222 79906 136500 79962
rect 136556 79906 136561 79962
rect 136222 79904 136561 79906
rect 134934 79792 135043 79797
rect 134934 79736 134982 79792
rect 135038 79736 135043 79792
rect 134934 79734 135043 79736
rect 134977 79731 135043 79734
rect 135294 79732 135300 79796
rect 135364 79794 135370 79796
rect 135440 79794 135500 79867
rect 135364 79734 135500 79794
rect 135364 79732 135370 79734
rect 134333 79658 134399 79661
rect 134152 79656 134399 79658
rect 134152 79600 134338 79656
rect 134394 79600 134399 79656
rect 134152 79598 134399 79600
rect 134750 79656 134859 79661
rect 134750 79600 134798 79656
rect 134854 79600 134859 79656
rect 134750 79598 134859 79600
rect 135670 79658 135730 79867
rect 136222 79794 136282 79904
rect 136495 79901 136561 79904
rect 136771 79962 136837 79967
rect 136771 79906 136776 79962
rect 136832 79906 136837 79962
rect 136771 79901 136837 79906
rect 136955 79962 137021 79967
rect 136955 79906 136960 79962
rect 137016 79906 137021 79962
rect 137415 79964 137481 79967
rect 139071 79964 139137 79967
rect 139439 79964 139505 79967
rect 140911 79964 140977 79967
rect 137415 79962 137754 79964
rect 137231 79930 137297 79933
rect 136955 79901 137021 79906
rect 137188 79928 137297 79930
rect 136449 79794 136515 79797
rect 136222 79792 136515 79794
rect 136222 79736 136454 79792
rect 136510 79736 136515 79792
rect 136222 79734 136515 79736
rect 136449 79731 136515 79734
rect 135805 79658 135871 79661
rect 135670 79656 135871 79658
rect 135670 79600 135810 79656
rect 135866 79600 135871 79656
rect 135670 79598 135871 79600
rect 134333 79595 134399 79598
rect 134793 79595 134859 79598
rect 135805 79595 135871 79598
rect 136633 79658 136699 79661
rect 136774 79658 136834 79901
rect 136958 79797 137018 79901
rect 137188 79872 137236 79928
rect 137292 79872 137297 79928
rect 137415 79906 137420 79962
rect 137476 79906 137754 79962
rect 139071 79962 139180 79964
rect 138059 79932 138125 79933
rect 138054 79930 138060 79932
rect 137415 79904 137754 79906
rect 137415 79901 137481 79904
rect 137188 79867 137297 79872
rect 136958 79792 137067 79797
rect 136958 79736 137006 79792
rect 137062 79736 137067 79792
rect 136958 79734 137067 79736
rect 137001 79731 137067 79734
rect 136633 79656 136834 79658
rect 136633 79600 136638 79656
rect 136694 79600 136834 79656
rect 136633 79598 136834 79600
rect 137188 79658 137248 79867
rect 137369 79658 137435 79661
rect 137188 79656 137435 79658
rect 137188 79600 137374 79656
rect 137430 79600 137435 79656
rect 137188 79598 137435 79600
rect 137694 79658 137754 79904
rect 137968 79870 138060 79930
rect 138054 79868 138060 79870
rect 138124 79868 138130 79932
rect 139071 79906 139076 79962
rect 139132 79932 139180 79962
rect 139439 79962 139686 79964
rect 139132 79906 139164 79932
rect 139071 79901 139164 79906
rect 139120 79870 139164 79901
rect 139158 79868 139164 79870
rect 139228 79868 139234 79932
rect 139439 79906 139444 79962
rect 139500 79906 139686 79962
rect 140911 79962 141020 79964
rect 139439 79904 139686 79906
rect 139439 79901 139505 79904
rect 138059 79867 138125 79868
rect 139347 79826 139413 79831
rect 137921 79796 137987 79797
rect 137870 79794 137876 79796
rect 137830 79734 137876 79794
rect 137940 79792 137987 79796
rect 137982 79736 137987 79792
rect 137870 79732 137876 79734
rect 137940 79732 137987 79736
rect 138974 79732 138980 79796
rect 139044 79794 139050 79796
rect 139347 79794 139352 79826
rect 139044 79770 139352 79794
rect 139408 79770 139413 79826
rect 139044 79765 139413 79770
rect 139626 79794 139686 79904
rect 140083 79894 140149 79899
rect 140083 79838 140088 79894
rect 140144 79838 140149 79894
rect 140630 79868 140636 79932
rect 140700 79930 140706 79932
rect 140911 79930 140916 79962
rect 140700 79906 140916 79930
rect 140972 79906 141020 79962
rect 141555 79962 141621 79967
rect 141279 79930 141345 79933
rect 140700 79870 141020 79906
rect 141236 79928 141345 79930
rect 141236 79872 141284 79928
rect 141340 79872 141345 79928
rect 141555 79906 141560 79962
rect 141616 79906 141621 79962
rect 142107 79962 142173 79967
rect 141555 79901 141621 79906
rect 141923 79930 141989 79933
rect 141923 79928 142032 79930
rect 140700 79868 140706 79870
rect 140083 79833 140149 79838
rect 141236 79867 141345 79872
rect 139945 79794 140011 79797
rect 139626 79792 140011 79794
rect 139044 79734 139410 79765
rect 139626 79736 139950 79792
rect 140006 79736 140011 79792
rect 139626 79734 140011 79736
rect 139044 79732 139050 79734
rect 137921 79731 137987 79732
rect 139945 79731 140011 79734
rect 140086 79661 140146 79833
rect 141236 79794 141296 79867
rect 141558 79797 141618 79901
rect 141923 79872 141928 79928
rect 141984 79872 142032 79928
rect 142107 79906 142112 79962
rect 142168 79906 142173 79962
rect 142107 79901 142173 79906
rect 142935 79962 143001 79967
rect 142935 79906 142940 79962
rect 142996 79906 143001 79962
rect 144131 79962 144197 79967
rect 142935 79901 143001 79906
rect 141923 79867 142032 79872
rect 141972 79797 142032 79867
rect 142475 79894 142541 79899
rect 142475 79838 142480 79894
rect 142536 79838 142541 79894
rect 143206 79868 143212 79932
rect 143276 79930 143282 79932
rect 143395 79930 143461 79933
rect 144131 79932 144136 79962
rect 144192 79932 144197 79962
rect 144683 79962 144749 79967
rect 143276 79928 143461 79930
rect 143276 79872 143400 79928
rect 143456 79872 143461 79928
rect 143276 79870 143461 79872
rect 143276 79868 143282 79870
rect 143395 79867 143461 79870
rect 144126 79868 144132 79932
rect 144196 79930 144202 79932
rect 144499 79930 144565 79933
rect 144683 79932 144688 79962
rect 144744 79932 144749 79962
rect 144196 79870 144254 79930
rect 144318 79928 144565 79930
rect 144318 79872 144504 79928
rect 144560 79872 144565 79928
rect 144318 79870 144565 79872
rect 144196 79868 144202 79870
rect 142475 79833 142541 79838
rect 141366 79794 141372 79796
rect 141236 79734 141372 79794
rect 141366 79732 141372 79734
rect 141436 79732 141442 79796
rect 141558 79792 141667 79797
rect 141558 79736 141606 79792
rect 141662 79736 141667 79792
rect 141558 79734 141667 79736
rect 141601 79731 141667 79734
rect 141969 79792 142035 79797
rect 141969 79736 141974 79792
rect 142030 79736 142035 79792
rect 141969 79731 142035 79736
rect 137921 79658 137987 79661
rect 137694 79656 137987 79658
rect 137694 79600 137926 79656
rect 137982 79600 137987 79656
rect 137694 79598 137987 79600
rect 136633 79595 136699 79598
rect 137369 79595 137435 79598
rect 137921 79595 137987 79598
rect 138606 79596 138612 79660
rect 138676 79658 138682 79660
rect 139025 79658 139091 79661
rect 139577 79660 139643 79661
rect 139526 79658 139532 79660
rect 138676 79656 139091 79658
rect 138676 79600 139030 79656
rect 139086 79600 139091 79656
rect 138676 79598 139091 79600
rect 139486 79598 139532 79658
rect 139596 79656 139643 79660
rect 139638 79600 139643 79656
rect 138676 79596 138682 79598
rect 139025 79595 139091 79598
rect 139526 79596 139532 79598
rect 139596 79596 139643 79600
rect 139577 79595 139643 79596
rect 140037 79656 140146 79661
rect 140037 79600 140042 79656
rect 140098 79600 140146 79656
rect 140037 79598 140146 79600
rect 140957 79658 141023 79661
rect 141417 79658 141483 79661
rect 140957 79656 141483 79658
rect 140957 79600 140962 79656
rect 141018 79600 141422 79656
rect 141478 79600 141483 79656
rect 140957 79598 141483 79600
rect 140037 79595 140103 79598
rect 140957 79595 141023 79598
rect 141417 79595 141483 79598
rect 142337 79658 142403 79661
rect 142478 79658 142538 79833
rect 142838 79732 142844 79796
rect 142908 79794 142914 79796
rect 143303 79794 143369 79797
rect 144318 79796 144378 79870
rect 144499 79867 144565 79870
rect 144678 79868 144684 79932
rect 144748 79930 144754 79932
rect 144748 79870 144806 79930
rect 144748 79868 144754 79870
rect 142908 79792 143369 79794
rect 142908 79736 143308 79792
rect 143364 79736 143369 79792
rect 142908 79734 143369 79736
rect 142908 79732 142914 79734
rect 143303 79731 143369 79734
rect 144310 79732 144316 79796
rect 144380 79732 144386 79796
rect 144494 79732 144500 79796
rect 144564 79794 144570 79796
rect 144870 79794 144930 80006
rect 145414 80004 145420 80006
rect 145484 80004 145490 80068
rect 148366 80066 148610 80100
rect 147998 80040 148610 80066
rect 147998 80006 148426 80040
rect 146339 79962 146405 79967
rect 145046 79868 145052 79932
rect 145116 79930 145122 79932
rect 145511 79930 145577 79933
rect 146063 79930 146129 79933
rect 145116 79928 145577 79930
rect 145116 79872 145516 79928
rect 145572 79872 145577 79928
rect 145116 79870 145577 79872
rect 145116 79868 145122 79870
rect 145511 79867 145577 79870
rect 145790 79928 146129 79930
rect 145790 79872 146068 79928
rect 146124 79872 146129 79928
rect 146339 79906 146344 79962
rect 146400 79906 146405 79962
rect 147351 79962 147417 79967
rect 146339 79901 146405 79906
rect 145790 79870 146129 79872
rect 145327 79794 145393 79797
rect 144564 79734 144930 79794
rect 145054 79792 145393 79794
rect 145054 79736 145332 79792
rect 145388 79736 145393 79792
rect 145054 79734 145393 79736
rect 144564 79732 144570 79734
rect 142337 79656 142538 79658
rect 142337 79600 142342 79656
rect 142398 79600 142538 79656
rect 142337 79598 142538 79600
rect 143809 79658 143875 79661
rect 144453 79658 144519 79661
rect 143809 79656 144519 79658
rect 143809 79600 143814 79656
rect 143870 79600 144458 79656
rect 144514 79600 144519 79656
rect 143809 79598 144519 79600
rect 145054 79658 145114 79734
rect 145327 79731 145393 79734
rect 145598 79732 145604 79796
rect 145668 79794 145674 79796
rect 145790 79794 145850 79870
rect 146063 79867 146129 79870
rect 145668 79734 145850 79794
rect 145668 79732 145674 79734
rect 146342 79661 146402 79901
rect 146523 79894 146589 79899
rect 146523 79838 146528 79894
rect 146584 79838 146589 79894
rect 147070 79868 147076 79932
rect 147140 79930 147146 79932
rect 147351 79930 147356 79962
rect 147140 79906 147356 79930
rect 147412 79906 147417 79962
rect 147140 79901 147417 79906
rect 147535 79962 147601 79967
rect 147535 79906 147540 79962
rect 147596 79906 147601 79962
rect 147535 79901 147601 79906
rect 147811 79962 147877 79967
rect 147811 79906 147816 79962
rect 147872 79906 147877 79962
rect 147811 79901 147877 79906
rect 147140 79870 147414 79901
rect 147140 79868 147146 79870
rect 146523 79833 146589 79838
rect 145281 79658 145347 79661
rect 145054 79656 145347 79658
rect 145054 79600 145286 79656
rect 145342 79600 145347 79656
rect 145054 79598 145347 79600
rect 142337 79595 142403 79598
rect 143809 79595 143875 79598
rect 144453 79595 144519 79598
rect 145281 79595 145347 79598
rect 145414 79596 145420 79660
rect 145484 79658 145490 79660
rect 145741 79658 145807 79661
rect 145484 79656 145807 79658
rect 145484 79600 145746 79656
rect 145802 79600 145807 79656
rect 145484 79598 145807 79600
rect 145484 79596 145490 79598
rect 145741 79595 145807 79598
rect 146293 79656 146402 79661
rect 146293 79600 146298 79656
rect 146354 79600 146402 79656
rect 146293 79598 146402 79600
rect 146526 79658 146586 79833
rect 147538 79797 147598 79901
rect 147814 79797 147874 79901
rect 147305 79796 147371 79797
rect 147254 79794 147260 79796
rect 147214 79734 147260 79794
rect 147324 79792 147371 79796
rect 147366 79736 147371 79792
rect 147254 79732 147260 79734
rect 147324 79732 147371 79736
rect 147538 79792 147647 79797
rect 147538 79736 147586 79792
rect 147642 79736 147647 79792
rect 147538 79734 147647 79736
rect 147814 79792 147923 79797
rect 147814 79736 147862 79792
rect 147918 79736 147923 79792
rect 147814 79734 147923 79736
rect 147305 79731 147371 79732
rect 147581 79731 147647 79734
rect 147857 79731 147923 79734
rect 147121 79658 147187 79661
rect 146526 79656 147187 79658
rect 146526 79600 147126 79656
rect 147182 79600 147187 79656
rect 146526 79598 147187 79600
rect 146293 79595 146359 79598
rect 147121 79595 147187 79598
rect 147765 79658 147831 79661
rect 147998 79658 148058 80006
rect 148550 79967 148610 80040
rect 152874 79967 152934 80142
rect 163446 80140 163452 80204
rect 163516 80202 163522 80204
rect 163516 80142 164158 80202
rect 163516 80140 163522 80142
rect 164098 79967 164158 80142
rect 164558 79967 164618 80278
rect 172278 80276 172284 80278
rect 172348 80276 172354 80340
rect 172094 80202 172100 80204
rect 168606 80142 172100 80202
rect 148547 79962 148613 79967
rect 148823 79964 148889 79967
rect 148174 79868 148180 79932
rect 148244 79930 148250 79932
rect 148363 79930 148429 79933
rect 148244 79928 148429 79930
rect 148244 79872 148368 79928
rect 148424 79872 148429 79928
rect 148547 79906 148552 79962
rect 148608 79906 148613 79962
rect 148780 79962 148889 79964
rect 148780 79932 148828 79962
rect 148547 79901 148613 79906
rect 148244 79870 148429 79872
rect 148244 79868 148250 79870
rect 148363 79867 148429 79870
rect 148726 79868 148732 79932
rect 148796 79906 148828 79932
rect 148884 79906 148889 79962
rect 148796 79901 148889 79906
rect 149467 79962 149533 79967
rect 150295 79964 150361 79967
rect 149467 79906 149472 79962
rect 149528 79906 149533 79962
rect 150252 79962 150361 79964
rect 149467 79901 149533 79906
rect 148796 79870 148840 79901
rect 148796 79868 148802 79870
rect 148542 79732 148548 79796
rect 148612 79794 148618 79796
rect 149007 79794 149073 79797
rect 148612 79792 149073 79794
rect 148612 79736 149012 79792
rect 149068 79736 149073 79792
rect 148612 79734 149073 79736
rect 148612 79732 148618 79734
rect 149007 79731 149073 79734
rect 147765 79656 148058 79658
rect 147765 79600 147770 79656
rect 147826 79600 148058 79656
rect 147765 79598 148058 79600
rect 148961 79658 149027 79661
rect 149470 79658 149530 79901
rect 149646 79868 149652 79932
rect 149716 79930 149722 79932
rect 150252 79930 150300 79962
rect 149716 79906 150300 79930
rect 150356 79906 150361 79962
rect 151491 79962 151557 79967
rect 149716 79901 150361 79906
rect 149716 79870 150312 79901
rect 149716 79868 149722 79870
rect 150566 79868 150572 79932
rect 150636 79930 150642 79932
rect 150847 79930 150913 79933
rect 150636 79928 150913 79930
rect 150636 79872 150852 79928
rect 150908 79872 150913 79928
rect 151491 79906 151496 79962
rect 151552 79906 151557 79962
rect 152871 79962 152937 79967
rect 151859 79932 151925 79933
rect 151854 79930 151860 79932
rect 151491 79901 151557 79906
rect 150636 79870 150913 79872
rect 150636 79868 150642 79870
rect 150847 79867 150913 79870
rect 150014 79732 150020 79796
rect 150084 79794 150090 79796
rect 150203 79794 150269 79797
rect 150084 79792 150269 79794
rect 150084 79736 150208 79792
rect 150264 79736 150269 79792
rect 150084 79734 150269 79736
rect 150084 79732 150090 79734
rect 150203 79731 150269 79734
rect 151353 79794 151419 79797
rect 151494 79794 151554 79901
rect 151768 79870 151860 79930
rect 151854 79868 151860 79870
rect 151924 79868 151930 79932
rect 152595 79928 152661 79933
rect 152595 79872 152600 79928
rect 152656 79872 152661 79928
rect 152871 79906 152876 79962
rect 152932 79906 152937 79962
rect 153147 79962 153213 79967
rect 156183 79964 156249 79967
rect 153147 79932 153152 79962
rect 153208 79932 153213 79962
rect 155910 79962 156249 79964
rect 152871 79901 152937 79906
rect 151859 79867 151925 79868
rect 152595 79867 152661 79872
rect 153142 79868 153148 79932
rect 153212 79930 153218 79932
rect 153212 79870 153270 79930
rect 153212 79868 153218 79870
rect 153878 79868 153884 79932
rect 153948 79930 153954 79932
rect 154527 79930 154593 79933
rect 155723 79932 155789 79933
rect 155718 79930 155724 79932
rect 153948 79928 154593 79930
rect 153948 79872 154532 79928
rect 154588 79872 154593 79928
rect 153948 79870 154593 79872
rect 155632 79870 155724 79930
rect 153948 79868 153954 79870
rect 154527 79867 154593 79870
rect 155718 79868 155724 79870
rect 155788 79868 155794 79932
rect 155910 79906 156188 79962
rect 156244 79906 156249 79962
rect 155910 79904 156249 79906
rect 155723 79867 155789 79868
rect 151353 79792 151554 79794
rect 151353 79736 151358 79792
rect 151414 79736 151554 79792
rect 151353 79734 151554 79736
rect 151675 79792 151741 79797
rect 151675 79736 151680 79792
rect 151736 79736 151741 79792
rect 151353 79731 151419 79734
rect 151675 79731 151741 79736
rect 148961 79656 149530 79658
rect 148961 79600 148966 79656
rect 149022 79600 149530 79656
rect 148961 79598 149530 79600
rect 147765 79595 147831 79598
rect 148961 79595 149027 79598
rect 151486 79596 151492 79660
rect 151556 79658 151562 79660
rect 151678 79658 151738 79731
rect 151556 79598 151738 79658
rect 152598 79658 152658 79867
rect 152774 79732 152780 79796
rect 152844 79794 152850 79796
rect 152917 79794 152983 79797
rect 152844 79792 152983 79794
rect 152844 79736 152922 79792
rect 152978 79736 152983 79792
rect 152844 79734 152983 79736
rect 152844 79732 152850 79734
rect 152917 79731 152983 79734
rect 153929 79794 153995 79797
rect 154481 79796 154547 79797
rect 154062 79794 154068 79796
rect 153929 79792 154068 79794
rect 153929 79736 153934 79792
rect 153990 79736 154068 79792
rect 153929 79734 154068 79736
rect 153929 79731 153995 79734
rect 154062 79732 154068 79734
rect 154132 79732 154138 79796
rect 154430 79794 154436 79796
rect 154390 79734 154436 79794
rect 154500 79792 154547 79796
rect 154542 79736 154547 79792
rect 154430 79732 154436 79734
rect 154500 79732 154547 79736
rect 154481 79731 154547 79732
rect 155910 79661 155970 79904
rect 156183 79901 156249 79904
rect 156367 79964 156433 79967
rect 156367 79962 156476 79964
rect 156367 79906 156372 79962
rect 156428 79906 156476 79962
rect 157103 79962 157169 79967
rect 156367 79901 156476 79906
rect 153101 79658 153167 79661
rect 152598 79656 153167 79658
rect 152598 79600 153106 79656
rect 153162 79600 153167 79656
rect 152598 79598 153167 79600
rect 151556 79596 151562 79598
rect 153101 79595 153167 79598
rect 154246 79596 154252 79660
rect 154316 79658 154322 79660
rect 154389 79658 154455 79661
rect 154316 79656 154455 79658
rect 154316 79600 154394 79656
rect 154450 79600 154455 79656
rect 154316 79598 154455 79600
rect 155910 79656 156019 79661
rect 155910 79600 155958 79656
rect 156014 79600 156019 79656
rect 155910 79598 156019 79600
rect 156416 79658 156476 79901
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157103 79930 157108 79962
rect 156892 79906 157108 79930
rect 157164 79906 157169 79962
rect 156892 79901 157169 79906
rect 157287 79964 157353 79967
rect 157287 79962 157396 79964
rect 157287 79906 157292 79962
rect 157348 79906 157396 79962
rect 158575 79962 158641 79967
rect 157287 79901 157396 79906
rect 156892 79870 157166 79901
rect 156892 79868 156898 79870
rect 156597 79658 156663 79661
rect 156416 79656 156663 79658
rect 156416 79600 156602 79656
rect 156658 79600 156663 79656
rect 156416 79598 156663 79600
rect 154316 79596 154322 79598
rect 154389 79595 154455 79598
rect 155953 79595 156019 79598
rect 156597 79595 156663 79598
rect 156822 79596 156828 79660
rect 156892 79658 156898 79660
rect 157336 79658 157396 79901
rect 157926 79868 157932 79932
rect 157996 79930 158002 79932
rect 158115 79930 158181 79933
rect 158299 79932 158365 79933
rect 157996 79928 158181 79930
rect 157996 79872 158120 79928
rect 158176 79872 158181 79928
rect 157996 79870 158181 79872
rect 157996 79868 158002 79870
rect 158115 79867 158181 79870
rect 158294 79868 158300 79932
rect 158364 79930 158370 79932
rect 158364 79870 158456 79930
rect 158575 79906 158580 79962
rect 158636 79906 158641 79962
rect 159771 79962 159837 79967
rect 159311 79930 159377 79933
rect 158575 79901 158641 79906
rect 159268 79928 159377 79930
rect 158364 79868 158370 79870
rect 158299 79867 158365 79868
rect 157563 79794 157629 79797
rect 157793 79794 157859 79797
rect 157563 79792 157859 79794
rect 157563 79736 157568 79792
rect 157624 79736 157798 79792
rect 157854 79736 157859 79792
rect 157563 79734 157859 79736
rect 157563 79731 157629 79734
rect 157793 79731 157859 79734
rect 158294 79732 158300 79796
rect 158364 79794 158370 79796
rect 158578 79794 158638 79901
rect 158943 79894 159009 79899
rect 158943 79838 158948 79894
rect 159004 79838 159009 79894
rect 158943 79833 159009 79838
rect 159268 79872 159316 79928
rect 159372 79872 159377 79928
rect 159268 79867 159377 79872
rect 159495 79928 159561 79933
rect 159495 79872 159500 79928
rect 159556 79872 159561 79928
rect 159771 79906 159776 79962
rect 159832 79906 159837 79962
rect 161427 79962 161493 79967
rect 159771 79901 159837 79906
rect 159495 79867 159561 79872
rect 158364 79734 158638 79794
rect 158364 79732 158370 79734
rect 156892 79598 157396 79658
rect 156892 79596 156898 79598
rect 157742 79596 157748 79660
rect 157812 79658 157818 79660
rect 157885 79658 157951 79661
rect 157812 79656 157951 79658
rect 157812 79600 157890 79656
rect 157946 79600 157951 79656
rect 157812 79598 157951 79600
rect 157812 79596 157818 79598
rect 157885 79595 157951 79598
rect 158713 79658 158779 79661
rect 158946 79658 159006 79833
rect 159268 79661 159328 79867
rect 159498 79661 159558 79867
rect 159774 79797 159834 79901
rect 159950 79868 159956 79932
rect 160020 79930 160026 79932
rect 160231 79930 160297 79933
rect 160875 79932 160941 79933
rect 161059 79932 161125 79933
rect 161427 79932 161432 79962
rect 161488 79932 161493 79962
rect 164095 79962 164161 79967
rect 160870 79930 160876 79932
rect 160020 79928 160297 79930
rect 160020 79872 160236 79928
rect 160292 79872 160297 79928
rect 160020 79870 160297 79872
rect 160784 79870 160876 79930
rect 160020 79868 160026 79870
rect 160231 79867 160297 79870
rect 160870 79868 160876 79870
rect 160940 79868 160946 79932
rect 161054 79868 161060 79932
rect 161124 79930 161130 79932
rect 161124 79870 161216 79930
rect 161124 79868 161130 79870
rect 161422 79868 161428 79932
rect 161492 79930 161498 79932
rect 161611 79930 161677 79933
rect 161790 79930 161796 79932
rect 161492 79870 161550 79930
rect 161611 79928 161796 79930
rect 161611 79872 161616 79928
rect 161672 79872 161796 79928
rect 161611 79870 161796 79872
rect 161492 79868 161498 79870
rect 160875 79867 160941 79868
rect 161059 79867 161125 79868
rect 161611 79867 161677 79870
rect 161790 79868 161796 79870
rect 161860 79868 161866 79932
rect 163727 79930 163793 79933
rect 163500 79928 163793 79930
rect 163500 79872 163732 79928
rect 163788 79872 163793 79928
rect 164095 79906 164100 79962
rect 164156 79906 164161 79962
rect 164095 79901 164161 79906
rect 164555 79962 164621 79967
rect 164555 79906 164560 79962
rect 164616 79906 164621 79962
rect 164555 79901 164621 79906
rect 164739 79962 164805 79967
rect 165015 79964 165081 79967
rect 164739 79906 164744 79962
rect 164800 79906 164805 79962
rect 164739 79901 164805 79906
rect 164880 79962 165081 79964
rect 164880 79906 165020 79962
rect 165076 79906 165081 79962
rect 167315 79962 167381 79967
rect 165475 79932 165541 79933
rect 166027 79932 166093 79933
rect 166211 79932 166277 79933
rect 165470 79930 165476 79932
rect 164880 79904 165081 79906
rect 163500 79870 163793 79872
rect 162439 79826 162505 79831
rect 159774 79792 159883 79797
rect 159774 79736 159822 79792
rect 159878 79736 159883 79792
rect 159774 79734 159883 79736
rect 159817 79731 159883 79734
rect 160502 79732 160508 79796
rect 160572 79794 160578 79796
rect 160921 79794 160987 79797
rect 160572 79792 160987 79794
rect 160572 79736 160926 79792
rect 160982 79736 160987 79792
rect 162439 79770 162444 79826
rect 162500 79794 162505 79826
rect 162710 79794 162716 79796
rect 162500 79770 162716 79794
rect 162439 79765 162716 79770
rect 160572 79734 160987 79736
rect 162442 79734 162716 79765
rect 160572 79732 160578 79734
rect 160921 79731 160987 79734
rect 162710 79732 162716 79734
rect 162780 79732 162786 79796
rect 162853 79794 162919 79797
rect 163078 79794 163084 79796
rect 162853 79792 163084 79794
rect 162853 79736 162858 79792
rect 162914 79736 163084 79792
rect 162853 79734 163084 79736
rect 162853 79731 162919 79734
rect 163078 79732 163084 79734
rect 163148 79732 163154 79796
rect 163500 79794 163560 79870
rect 163727 79867 163793 79870
rect 163681 79794 163747 79797
rect 163500 79792 163747 79794
rect 163500 79736 163686 79792
rect 163742 79736 163747 79792
rect 163500 79734 163747 79736
rect 163681 79731 163747 79734
rect 164742 79661 164802 79901
rect 164880 79794 164940 79904
rect 165015 79901 165081 79904
rect 165384 79870 165476 79930
rect 165470 79868 165476 79870
rect 165540 79868 165546 79932
rect 166022 79930 166028 79932
rect 165936 79870 166028 79930
rect 166022 79868 166028 79870
rect 166092 79868 166098 79932
rect 166206 79868 166212 79932
rect 166276 79930 166282 79932
rect 166276 79870 166368 79930
rect 166947 79928 167013 79933
rect 167315 79932 167320 79962
rect 167376 79932 167381 79962
rect 166947 79872 166952 79928
rect 167008 79872 167013 79928
rect 166276 79868 166282 79870
rect 165475 79867 165541 79868
rect 166027 79867 166093 79868
rect 166211 79867 166277 79868
rect 166947 79867 167013 79872
rect 167310 79868 167316 79932
rect 167380 79930 167386 79932
rect 167380 79870 167438 79930
rect 167380 79868 167386 79870
rect 168046 79868 168052 79932
rect 168116 79930 168122 79932
rect 168235 79930 168301 79933
rect 168116 79928 168301 79930
rect 168116 79872 168240 79928
rect 168296 79872 168301 79928
rect 168116 79870 168301 79872
rect 168116 79868 168122 79870
rect 168235 79867 168301 79870
rect 164880 79734 165170 79794
rect 165110 79661 165170 79734
rect 166390 79732 166396 79796
rect 166460 79794 166466 79796
rect 166950 79794 167010 79867
rect 166460 79734 167010 79794
rect 166460 79732 166466 79734
rect 167678 79732 167684 79796
rect 167748 79794 167754 79796
rect 168005 79794 168071 79797
rect 167748 79792 168071 79794
rect 167748 79736 168010 79792
rect 168066 79736 168071 79792
rect 167748 79734 168071 79736
rect 167748 79732 167754 79734
rect 168005 79731 168071 79734
rect 168373 79794 168439 79797
rect 168606 79794 168666 80142
rect 172094 80140 172100 80142
rect 172164 80140 172170 80204
rect 173014 80202 173020 80204
rect 172240 80142 173020 80202
rect 172240 79967 172300 80142
rect 173014 80140 173020 80142
rect 173084 80140 173090 80204
rect 168787 79962 168853 79967
rect 168787 79906 168792 79962
rect 168848 79906 168853 79962
rect 168787 79901 168853 79906
rect 168971 79962 169037 79967
rect 168971 79906 168976 79962
rect 169032 79930 169037 79962
rect 170443 79962 170509 79967
rect 169891 79932 169957 79933
rect 169886 79930 169892 79932
rect 169032 79906 169724 79930
rect 168971 79901 169724 79906
rect 168373 79792 168666 79794
rect 168373 79736 168378 79792
rect 168434 79736 168666 79792
rect 168373 79734 168666 79736
rect 168373 79731 168439 79734
rect 168790 79661 168850 79901
rect 168974 79870 169724 79901
rect 169800 79870 169892 79930
rect 169431 79794 169497 79797
rect 158713 79656 159006 79658
rect 158713 79600 158718 79656
rect 158774 79600 159006 79656
rect 158713 79598 159006 79600
rect 159265 79656 159331 79661
rect 159265 79600 159270 79656
rect 159326 79600 159331 79656
rect 158713 79595 158779 79598
rect 159265 79595 159331 79600
rect 159449 79656 159558 79661
rect 159449 79600 159454 79656
rect 159510 79600 159558 79656
rect 159449 79598 159558 79600
rect 160093 79658 160159 79661
rect 160318 79658 160324 79660
rect 160093 79656 160324 79658
rect 160093 79600 160098 79656
rect 160154 79600 160324 79656
rect 160093 79598 160324 79600
rect 159449 79595 159515 79598
rect 160093 79595 160159 79598
rect 160318 79596 160324 79598
rect 160388 79596 160394 79660
rect 160686 79596 160692 79660
rect 160756 79658 160762 79660
rect 161105 79658 161171 79661
rect 160756 79656 161171 79658
rect 160756 79600 161110 79656
rect 161166 79600 161171 79656
rect 160756 79598 161171 79600
rect 160756 79596 160762 79598
rect 161105 79595 161171 79598
rect 162526 79596 162532 79660
rect 162596 79658 162602 79660
rect 162669 79658 162735 79661
rect 162596 79656 162735 79658
rect 162596 79600 162674 79656
rect 162730 79600 162735 79656
rect 162596 79598 162735 79600
rect 162596 79596 162602 79598
rect 162669 79595 162735 79598
rect 163262 79596 163268 79660
rect 163332 79658 163338 79660
rect 163497 79658 163563 79661
rect 163332 79656 163563 79658
rect 163332 79600 163502 79656
rect 163558 79600 163563 79656
rect 163332 79598 163563 79600
rect 163332 79596 163338 79598
rect 163497 79595 163563 79598
rect 163630 79596 163636 79660
rect 163700 79658 163706 79660
rect 164049 79658 164115 79661
rect 163700 79656 164115 79658
rect 163700 79600 164054 79656
rect 164110 79600 164115 79656
rect 163700 79598 164115 79600
rect 164742 79656 164851 79661
rect 164742 79600 164790 79656
rect 164846 79600 164851 79656
rect 164742 79598 164851 79600
rect 163700 79596 163706 79598
rect 164049 79595 164115 79598
rect 164785 79595 164851 79598
rect 165061 79656 165170 79661
rect 165061 79600 165066 79656
rect 165122 79600 165170 79656
rect 165061 79598 165170 79600
rect 165061 79595 165127 79598
rect 166574 79596 166580 79660
rect 166644 79658 166650 79660
rect 166901 79658 166967 79661
rect 166644 79656 166967 79658
rect 166644 79600 166906 79656
rect 166962 79600 166967 79656
rect 166644 79598 166967 79600
rect 166644 79596 166650 79598
rect 166901 79595 166967 79598
rect 168741 79656 168850 79661
rect 168741 79600 168746 79656
rect 168802 79600 168850 79656
rect 168741 79598 168850 79600
rect 169204 79792 169497 79794
rect 169204 79736 169436 79792
rect 169492 79736 169497 79792
rect 169204 79734 169497 79736
rect 169664 79794 169724 79870
rect 169886 79868 169892 79870
rect 169956 79868 169962 79932
rect 170443 79906 170448 79962
rect 170504 79930 170509 79962
rect 171363 79962 171429 79967
rect 170806 79930 170812 79932
rect 170504 79906 170812 79930
rect 170443 79901 170812 79906
rect 170446 79870 170812 79901
rect 170806 79868 170812 79870
rect 170876 79868 170882 79932
rect 171087 79928 171153 79933
rect 171363 79932 171368 79962
rect 171424 79932 171429 79962
rect 172191 79962 172300 79967
rect 171087 79872 171092 79928
rect 171148 79872 171153 79928
rect 169891 79867 169957 79868
rect 171087 79867 171153 79872
rect 171358 79868 171364 79932
rect 171428 79930 171434 79932
rect 171547 79930 171613 79933
rect 171910 79930 171916 79932
rect 171428 79870 171486 79930
rect 171547 79928 171916 79930
rect 171547 79872 171552 79928
rect 171608 79872 171916 79928
rect 171547 79870 171916 79872
rect 171428 79868 171434 79870
rect 171547 79867 171613 79870
rect 171910 79868 171916 79870
rect 171980 79868 171986 79932
rect 172191 79906 172196 79962
rect 172252 79906 172300 79962
rect 172191 79904 172300 79906
rect 172375 79930 172441 79933
rect 173019 79932 173085 79933
rect 172646 79930 172652 79932
rect 172375 79928 172652 79930
rect 172191 79901 172257 79904
rect 172375 79872 172380 79928
rect 172436 79872 172652 79928
rect 172375 79870 172652 79872
rect 172375 79867 172441 79870
rect 172646 79868 172652 79870
rect 172716 79868 172722 79932
rect 173014 79930 173020 79932
rect 172928 79870 173020 79930
rect 173014 79868 173020 79870
rect 173084 79868 173090 79932
rect 173019 79867 173085 79868
rect 169845 79794 169911 79797
rect 169664 79792 169911 79794
rect 169664 79736 169850 79792
rect 169906 79736 169911 79792
rect 169664 79734 169911 79736
rect 169204 79658 169264 79734
rect 169431 79731 169497 79734
rect 169845 79731 169911 79734
rect 170622 79732 170628 79796
rect 170692 79794 170698 79796
rect 170811 79794 170877 79797
rect 170692 79792 170877 79794
rect 170692 79736 170816 79792
rect 170872 79736 170877 79792
rect 170692 79734 170877 79736
rect 171090 79794 171150 79867
rect 172646 79794 172652 79796
rect 171090 79734 172652 79794
rect 170692 79732 170698 79734
rect 170811 79731 170877 79734
rect 172646 79732 172652 79734
rect 172716 79732 172722 79796
rect 172973 79794 173039 79797
rect 173160 79794 173220 80414
rect 173295 79964 173361 79967
rect 173295 79962 173404 79964
rect 173295 79906 173300 79962
rect 173356 79932 173404 79962
rect 173939 79932 174005 79933
rect 173356 79906 173388 79932
rect 173295 79901 173388 79906
rect 173344 79870 173388 79901
rect 173382 79868 173388 79870
rect 173452 79868 173458 79932
rect 173934 79930 173940 79932
rect 173848 79870 173940 79930
rect 173934 79868 173940 79870
rect 174004 79868 174010 79932
rect 173939 79867 174005 79868
rect 172973 79792 173220 79794
rect 172973 79736 172978 79792
rect 173034 79736 173220 79792
rect 172973 79734 173220 79736
rect 172973 79731 173039 79734
rect 173566 79732 173572 79796
rect 173636 79794 173642 79796
rect 173985 79794 174051 79797
rect 173636 79792 174051 79794
rect 173636 79736 173990 79792
rect 174046 79736 174051 79792
rect 173636 79734 174051 79736
rect 173636 79732 173642 79734
rect 173985 79731 174051 79734
rect 169385 79658 169451 79661
rect 169204 79656 169451 79658
rect 169204 79600 169390 79656
rect 169446 79600 169451 79656
rect 169204 79598 169451 79600
rect 168741 79595 168807 79598
rect 169385 79595 169451 79598
rect 169518 79596 169524 79660
rect 169588 79658 169594 79660
rect 169661 79658 169727 79661
rect 169588 79656 169727 79658
rect 169588 79600 169666 79656
rect 169722 79600 169727 79656
rect 169588 79598 169727 79600
rect 169588 79596 169594 79598
rect 169661 79595 169727 79598
rect 171133 79658 171199 79661
rect 174353 79658 174419 79661
rect 171133 79656 174419 79658
rect 171133 79600 171138 79656
rect 171194 79600 174358 79656
rect 174414 79600 174419 79656
rect 171133 79598 174419 79600
rect 171133 79595 171199 79598
rect 174353 79595 174419 79598
rect 6913 79522 6979 79525
rect 168097 79522 168163 79525
rect 6913 79520 168163 79522
rect 6913 79464 6918 79520
rect 6974 79464 168102 79520
rect 168158 79464 168163 79520
rect 6913 79462 168163 79464
rect 6913 79459 6979 79462
rect 168097 79459 168163 79462
rect 171910 79460 171916 79524
rect 171980 79522 171986 79524
rect 172513 79522 172579 79525
rect 171980 79520 172579 79522
rect 171980 79464 172518 79520
rect 172574 79464 172579 79520
rect 171980 79462 172579 79464
rect 171980 79460 171986 79462
rect 172513 79459 172579 79462
rect 172646 79460 172652 79524
rect 172716 79522 172722 79524
rect 180425 79522 180491 79525
rect 172716 79520 180491 79522
rect 172716 79464 180430 79520
rect 180486 79464 180491 79520
rect 172716 79462 180491 79464
rect 172716 79460 172722 79462
rect 180425 79459 180491 79462
rect 3969 79386 4035 79389
rect 173525 79386 173591 79389
rect 3969 79384 173591 79386
rect 3969 79328 3974 79384
rect 4030 79328 173530 79384
rect 173586 79328 173591 79384
rect 3969 79326 173591 79328
rect 3969 79323 4035 79326
rect 173525 79323 173591 79326
rect 176285 79386 176351 79389
rect 580809 79386 580875 79389
rect 176285 79384 580875 79386
rect 176285 79328 176290 79384
rect 176346 79328 580814 79384
rect 580870 79328 580875 79384
rect 176285 79326 580875 79328
rect 176285 79323 176351 79326
rect 580809 79323 580875 79326
rect 3785 79250 3851 79253
rect 173382 79250 173388 79252
rect 3785 79248 173388 79250
rect 3785 79192 3790 79248
rect 3846 79192 173388 79248
rect 3785 79190 173388 79192
rect 3785 79187 3851 79190
rect 173382 79188 173388 79190
rect 173452 79188 173458 79252
rect 3601 79114 3667 79117
rect 171777 79114 171843 79117
rect 176101 79114 176167 79117
rect 3601 79112 171843 79114
rect 3601 79056 3606 79112
rect 3662 79056 171782 79112
rect 171838 79056 171843 79112
rect 3601 79054 171843 79056
rect 3601 79051 3667 79054
rect 171777 79051 171843 79054
rect 172102 79112 176167 79114
rect 172102 79056 176106 79112
rect 176162 79056 176167 79112
rect 172102 79054 176167 79056
rect 3417 78978 3483 78981
rect 171501 78978 171567 78981
rect 172102 78978 172162 79054
rect 176101 79051 176167 79054
rect 3417 78976 168666 78978
rect 3417 78920 3422 78976
rect 3478 78920 168666 78976
rect 3417 78918 168666 78920
rect 3417 78915 3483 78918
rect 128353 78842 128419 78845
rect 128854 78842 128860 78844
rect 128353 78840 128860 78842
rect 128353 78784 128358 78840
rect 128414 78784 128860 78840
rect 128353 78782 128860 78784
rect 128353 78779 128419 78782
rect 128854 78780 128860 78782
rect 128924 78780 128930 78844
rect 129733 78842 129799 78845
rect 130142 78842 130148 78844
rect 129733 78840 130148 78842
rect 129733 78784 129738 78840
rect 129794 78784 130148 78840
rect 129733 78782 130148 78784
rect 129733 78779 129799 78782
rect 130142 78780 130148 78782
rect 130212 78780 130218 78844
rect 136398 78780 136404 78844
rect 136468 78842 136474 78844
rect 136817 78842 136883 78845
rect 136468 78840 136883 78842
rect 136468 78784 136822 78840
rect 136878 78784 136883 78840
rect 136468 78782 136883 78784
rect 136468 78780 136474 78782
rect 136817 78779 136883 78782
rect 137686 78780 137692 78844
rect 137756 78842 137762 78844
rect 138105 78842 138171 78845
rect 137756 78840 138171 78842
rect 137756 78784 138110 78840
rect 138166 78784 138171 78840
rect 137756 78782 138171 78784
rect 137756 78780 137762 78782
rect 138105 78779 138171 78782
rect 140446 78780 140452 78844
rect 140516 78842 140522 78844
rect 140865 78842 140931 78845
rect 140516 78840 140931 78842
rect 140516 78784 140870 78840
rect 140926 78784 140931 78840
rect 140516 78782 140931 78784
rect 140516 78780 140522 78782
rect 140865 78779 140931 78782
rect 151302 78780 151308 78844
rect 151372 78842 151378 78844
rect 151721 78842 151787 78845
rect 151372 78840 151787 78842
rect 151372 78784 151726 78840
rect 151782 78784 151787 78840
rect 151372 78782 151787 78784
rect 151372 78780 151378 78782
rect 151721 78779 151787 78782
rect 159950 78780 159956 78844
rect 160020 78842 160026 78844
rect 160277 78842 160343 78845
rect 160020 78840 160343 78842
rect 160020 78784 160282 78840
rect 160338 78784 160343 78840
rect 160020 78782 160343 78784
rect 160020 78780 160026 78782
rect 160277 78779 160343 78782
rect 165102 78780 165108 78844
rect 165172 78842 165178 78844
rect 165521 78842 165587 78845
rect 165172 78840 165587 78842
rect 165172 78784 165526 78840
rect 165582 78784 165587 78840
rect 165172 78782 165587 78784
rect 168606 78842 168666 78918
rect 171501 78976 172162 78978
rect 171501 78920 171506 78976
rect 171562 78920 172162 78976
rect 171501 78918 172162 78920
rect 172237 78978 172303 78981
rect 173709 78978 173775 78981
rect 172237 78976 173775 78978
rect 172237 78920 172242 78976
rect 172298 78920 173714 78976
rect 173770 78920 173775 78976
rect 172237 78918 173775 78920
rect 171501 78915 171567 78918
rect 172237 78915 172303 78918
rect 173709 78915 173775 78918
rect 172697 78842 172763 78845
rect 168606 78840 172763 78842
rect 168606 78784 172702 78840
rect 172758 78784 172763 78840
rect 168606 78782 172763 78784
rect 165172 78780 165178 78782
rect 165521 78779 165587 78782
rect 172697 78779 172763 78782
rect 172830 78780 172836 78844
rect 172900 78842 172906 78844
rect 175917 78842 175983 78845
rect 397453 78842 397519 78845
rect 172900 78782 175842 78842
rect 172900 78780 172906 78782
rect 129222 78644 129228 78708
rect 129292 78706 129298 78708
rect 129365 78706 129431 78709
rect 130009 78708 130075 78709
rect 129958 78706 129964 78708
rect 129292 78704 129431 78706
rect 129292 78648 129370 78704
rect 129426 78648 129431 78704
rect 129292 78646 129431 78648
rect 129918 78646 129964 78706
rect 130028 78704 130075 78708
rect 130070 78648 130075 78704
rect 129292 78644 129298 78646
rect 129365 78643 129431 78646
rect 129958 78644 129964 78646
rect 130028 78644 130075 78648
rect 130009 78643 130075 78644
rect 131205 78706 131271 78709
rect 134057 78708 134123 78709
rect 131430 78706 131436 78708
rect 131205 78704 131436 78706
rect 131205 78648 131210 78704
rect 131266 78648 131436 78704
rect 131205 78646 131436 78648
rect 131205 78643 131271 78646
rect 131430 78644 131436 78646
rect 131500 78644 131506 78708
rect 134006 78706 134012 78708
rect 133966 78646 134012 78706
rect 134076 78704 134123 78708
rect 138013 78708 138079 78709
rect 138013 78706 138060 78708
rect 134118 78648 134123 78704
rect 134006 78644 134012 78646
rect 134076 78644 134123 78648
rect 137968 78704 138060 78706
rect 137968 78648 138018 78704
rect 137968 78646 138060 78648
rect 134057 78643 134123 78644
rect 138013 78644 138060 78646
rect 138124 78644 138130 78708
rect 138790 78644 138796 78708
rect 138860 78706 138866 78708
rect 139117 78706 139183 78709
rect 138860 78704 139183 78706
rect 138860 78648 139122 78704
rect 139178 78648 139183 78704
rect 138860 78646 139183 78648
rect 138860 78644 138866 78646
rect 138013 78643 138079 78644
rect 139117 78643 139183 78646
rect 151537 78706 151603 78709
rect 151905 78708 151971 78709
rect 151670 78706 151676 78708
rect 151537 78704 151676 78706
rect 151537 78648 151542 78704
rect 151598 78648 151676 78704
rect 151537 78646 151676 78648
rect 151537 78643 151603 78646
rect 151670 78644 151676 78646
rect 151740 78644 151746 78708
rect 151854 78644 151860 78708
rect 151924 78706 151971 78708
rect 151924 78704 152016 78706
rect 151966 78648 152016 78704
rect 151924 78646 152016 78648
rect 151924 78644 151971 78646
rect 156638 78644 156644 78708
rect 156708 78706 156714 78708
rect 156965 78706 157031 78709
rect 156708 78704 157031 78706
rect 156708 78648 156970 78704
rect 157026 78648 157031 78704
rect 156708 78646 157031 78648
rect 156708 78644 156714 78646
rect 151905 78643 151971 78644
rect 156965 78643 157031 78646
rect 160318 78644 160324 78708
rect 160388 78706 160394 78708
rect 160737 78706 160803 78709
rect 160388 78704 160803 78706
rect 160388 78648 160742 78704
rect 160798 78648 160803 78704
rect 160388 78646 160803 78648
rect 160388 78644 160394 78646
rect 160737 78643 160803 78646
rect 163262 78644 163268 78708
rect 163332 78706 163338 78708
rect 163405 78706 163471 78709
rect 163332 78704 163471 78706
rect 163332 78648 163410 78704
rect 163466 78648 163471 78704
rect 163332 78646 163471 78648
rect 163332 78644 163338 78646
rect 163405 78643 163471 78646
rect 168097 78706 168163 78709
rect 173014 78706 173020 78708
rect 168097 78704 173020 78706
rect 168097 78648 168102 78704
rect 168158 78648 173020 78704
rect 168097 78646 173020 78648
rect 168097 78643 168163 78646
rect 173014 78644 173020 78646
rect 173084 78644 173090 78708
rect 173198 78644 173204 78708
rect 173268 78706 173274 78708
rect 175641 78706 175707 78709
rect 173268 78704 175707 78706
rect 173268 78648 175646 78704
rect 175702 78648 175707 78704
rect 173268 78646 175707 78648
rect 175782 78706 175842 78782
rect 175917 78840 397519 78842
rect 175917 78784 175922 78840
rect 175978 78784 397458 78840
rect 397514 78784 397519 78840
rect 175917 78782 397519 78784
rect 175917 78779 175983 78782
rect 397453 78779 397519 78782
rect 462313 78706 462379 78709
rect 175782 78704 462379 78706
rect 175782 78648 462318 78704
rect 462374 78648 462379 78704
rect 175782 78646 462379 78648
rect 173268 78644 173274 78646
rect 175641 78643 175707 78646
rect 462313 78643 462379 78646
rect 44817 78570 44883 78573
rect 173566 78570 173572 78572
rect 44817 78568 173572 78570
rect 44817 78512 44822 78568
rect 44878 78512 173572 78568
rect 44817 78510 173572 78512
rect 44817 78507 44883 78510
rect 173566 78508 173572 78510
rect 173636 78508 173642 78572
rect 173934 78434 173940 78436
rect 128310 78374 173940 78434
rect 122097 78162 122163 78165
rect 127341 78162 127407 78165
rect 122097 78160 127407 78162
rect 122097 78104 122102 78160
rect 122158 78104 127346 78160
rect 127402 78104 127407 78160
rect 122097 78102 127407 78104
rect 122097 78099 122163 78102
rect 127341 78099 127407 78102
rect 119337 78026 119403 78029
rect 128310 78026 128370 78374
rect 173934 78372 173940 78374
rect 174004 78372 174010 78436
rect 133638 78236 133644 78300
rect 133708 78298 133714 78300
rect 140630 78298 140636 78300
rect 133708 78238 140636 78298
rect 133708 78236 133714 78238
rect 140630 78236 140636 78238
rect 140700 78236 140706 78300
rect 162945 78298 163011 78301
rect 171133 78298 171199 78301
rect 162945 78296 171199 78298
rect 162945 78240 162950 78296
rect 163006 78240 171138 78296
rect 171194 78240 171199 78296
rect 162945 78238 171199 78240
rect 162945 78235 163011 78238
rect 171133 78235 171199 78238
rect 171777 78298 171843 78301
rect 173157 78298 173223 78301
rect 171777 78296 173223 78298
rect 171777 78240 171782 78296
rect 171838 78240 173162 78296
rect 173218 78240 173223 78296
rect 171777 78238 173223 78240
rect 171777 78235 171843 78238
rect 173157 78235 173223 78238
rect 131665 78162 131731 78165
rect 132166 78162 132172 78164
rect 131665 78160 132172 78162
rect 131665 78104 131670 78160
rect 131726 78104 132172 78160
rect 131665 78102 132172 78104
rect 131665 78099 131731 78102
rect 132166 78100 132172 78102
rect 132236 78100 132242 78164
rect 141366 78100 141372 78164
rect 141436 78162 141442 78164
rect 141601 78162 141667 78165
rect 141436 78160 141667 78162
rect 141436 78104 141606 78160
rect 141662 78104 141667 78160
rect 141436 78102 141667 78104
rect 141436 78100 141442 78102
rect 141601 78099 141667 78102
rect 149830 78100 149836 78164
rect 149900 78162 149906 78164
rect 149973 78162 150039 78165
rect 150525 78164 150591 78165
rect 150525 78162 150572 78164
rect 149900 78160 150039 78162
rect 149900 78104 149978 78160
rect 150034 78104 150039 78160
rect 149900 78102 150039 78104
rect 150480 78160 150572 78162
rect 150480 78104 150530 78160
rect 150480 78102 150572 78104
rect 149900 78100 149906 78102
rect 149973 78099 150039 78102
rect 150525 78100 150572 78102
rect 150636 78100 150642 78164
rect 161289 78162 161355 78165
rect 255957 78162 256023 78165
rect 161289 78160 256023 78162
rect 161289 78104 161294 78160
rect 161350 78104 255962 78160
rect 256018 78104 256023 78160
rect 161289 78102 256023 78104
rect 150525 78099 150591 78100
rect 161289 78099 161355 78102
rect 255957 78099 256023 78102
rect 119337 78024 128370 78026
rect 119337 77968 119342 78024
rect 119398 77968 128370 78024
rect 119337 77966 128370 77968
rect 132585 78026 132651 78029
rect 133270 78026 133276 78028
rect 132585 78024 133276 78026
rect 132585 77968 132590 78024
rect 132646 77968 133276 78024
rect 132585 77966 133276 77968
rect 119337 77963 119403 77966
rect 132585 77963 132651 77966
rect 133270 77964 133276 77966
rect 133340 77964 133346 78028
rect 133965 78026 134031 78029
rect 134190 78026 134196 78028
rect 133965 78024 134196 78026
rect 133965 77968 133970 78024
rect 134026 77968 134196 78024
rect 133965 77966 134196 77968
rect 133965 77963 134031 77966
rect 134190 77964 134196 77966
rect 134260 77964 134266 78028
rect 134926 77964 134932 78028
rect 134996 78026 135002 78028
rect 171133 78026 171199 78029
rect 436737 78026 436803 78029
rect 134996 77966 138306 78026
rect 134996 77964 135002 77966
rect 10317 77890 10383 77893
rect 125041 77890 125107 77893
rect 10317 77888 125107 77890
rect 10317 77832 10322 77888
rect 10378 77832 125046 77888
rect 125102 77832 125107 77888
rect 10317 77830 125107 77832
rect 10317 77827 10383 77830
rect 125041 77827 125107 77830
rect 125501 77890 125567 77893
rect 125910 77890 125916 77892
rect 125501 77888 125916 77890
rect 125501 77832 125506 77888
rect 125562 77832 125916 77888
rect 125501 77830 125916 77832
rect 125501 77827 125567 77830
rect 125910 77828 125916 77830
rect 125980 77828 125986 77892
rect 127433 77890 127499 77893
rect 127566 77890 127572 77892
rect 127433 77888 127572 77890
rect 127433 77832 127438 77888
rect 127494 77832 127572 77888
rect 127433 77830 127572 77832
rect 127433 77827 127499 77830
rect 127566 77828 127572 77830
rect 127636 77828 127642 77892
rect 129733 77890 129799 77893
rect 133454 77890 133460 77892
rect 129733 77888 133460 77890
rect 129733 77832 129738 77888
rect 129794 77832 133460 77888
rect 129733 77830 133460 77832
rect 129733 77827 129799 77830
rect 133454 77828 133460 77830
rect 133524 77828 133530 77892
rect 136030 77828 136036 77892
rect 136100 77890 136106 77892
rect 138054 77890 138060 77892
rect 136100 77830 138060 77890
rect 136100 77828 136106 77830
rect 138054 77828 138060 77830
rect 138124 77828 138130 77892
rect 138246 77890 138306 77966
rect 171133 78024 436803 78026
rect 171133 77968 171138 78024
rect 171194 77968 436742 78024
rect 436798 77968 436803 78024
rect 171133 77966 436803 77968
rect 171133 77963 171199 77966
rect 436737 77963 436803 77966
rect 144545 77890 144611 77893
rect 138246 77888 144611 77890
rect 138246 77832 144550 77888
rect 144606 77832 144611 77888
rect 138246 77830 144611 77832
rect 144545 77827 144611 77830
rect 157926 77828 157932 77892
rect 157996 77890 158002 77892
rect 159173 77890 159239 77893
rect 157996 77888 159239 77890
rect 157996 77832 159178 77888
rect 159234 77832 159239 77888
rect 157996 77830 159239 77832
rect 157996 77828 158002 77830
rect 159173 77827 159239 77830
rect 162669 77890 162735 77893
rect 483013 77890 483079 77893
rect 162669 77888 483079 77890
rect 162669 77832 162674 77888
rect 162730 77832 483018 77888
rect 483074 77832 483079 77888
rect 162669 77830 483079 77832
rect 162669 77827 162735 77830
rect 483013 77827 483079 77830
rect 125777 77754 125843 77757
rect 126278 77754 126284 77756
rect 125777 77752 126284 77754
rect 125777 77696 125782 77752
rect 125838 77696 126284 77752
rect 125777 77694 126284 77696
rect 125777 77691 125843 77694
rect 126278 77692 126284 77694
rect 126348 77692 126354 77756
rect 131982 77692 131988 77756
rect 132052 77754 132058 77756
rect 142889 77754 142955 77757
rect 132052 77752 142955 77754
rect 132052 77696 142894 77752
rect 142950 77696 142955 77752
rect 132052 77694 142955 77696
rect 132052 77692 132058 77694
rect 142889 77691 142955 77694
rect 171685 77754 171751 77757
rect 174537 77754 174603 77757
rect 171685 77752 174603 77754
rect 171685 77696 171690 77752
rect 171746 77696 174542 77752
rect 174598 77696 174603 77752
rect 171685 77694 174603 77696
rect 171685 77691 171751 77694
rect 174537 77691 174603 77694
rect 168046 77420 168052 77484
rect 168116 77482 168122 77484
rect 168189 77482 168255 77485
rect 169937 77484 170003 77485
rect 170489 77484 170555 77485
rect 168116 77480 168255 77482
rect 168116 77424 168194 77480
rect 168250 77424 168255 77480
rect 168116 77422 168255 77424
rect 168116 77420 168122 77422
rect 168189 77419 168255 77422
rect 169886 77420 169892 77484
rect 169956 77482 170003 77484
rect 170438 77482 170444 77484
rect 169956 77480 170048 77482
rect 169998 77424 170048 77480
rect 169956 77422 170048 77424
rect 170398 77422 170444 77482
rect 170508 77480 170555 77484
rect 170550 77424 170555 77480
rect 169956 77420 170003 77422
rect 170438 77420 170444 77422
rect 170508 77420 170555 77424
rect 169937 77419 170003 77420
rect 170489 77419 170555 77420
rect 138054 77284 138060 77348
rect 138124 77346 138130 77348
rect 138124 77286 138490 77346
rect 138124 77284 138130 77286
rect 138430 77210 138490 77286
rect 149462 77284 149468 77348
rect 149532 77346 149538 77348
rect 150065 77346 150131 77349
rect 149532 77344 150131 77346
rect 149532 77288 150070 77344
rect 150126 77288 150131 77344
rect 149532 77286 150131 77288
rect 149532 77284 149538 77286
rect 150065 77283 150131 77286
rect 152590 77284 152596 77348
rect 152660 77346 152666 77348
rect 152917 77346 152983 77349
rect 157793 77348 157859 77349
rect 152660 77344 152983 77346
rect 152660 77288 152922 77344
rect 152978 77288 152983 77344
rect 152660 77286 152983 77288
rect 152660 77284 152666 77286
rect 152917 77283 152983 77286
rect 157742 77284 157748 77348
rect 157812 77346 157859 77348
rect 157812 77344 157904 77346
rect 157854 77288 157904 77344
rect 157812 77286 157904 77288
rect 157812 77284 157859 77286
rect 163078 77284 163084 77348
rect 163148 77346 163154 77348
rect 165613 77346 165679 77349
rect 163148 77344 165679 77346
rect 163148 77288 165618 77344
rect 165674 77288 165679 77344
rect 163148 77286 165679 77288
rect 163148 77284 163154 77286
rect 157793 77283 157859 77284
rect 165613 77283 165679 77286
rect 170397 77346 170463 77349
rect 170806 77346 170812 77348
rect 170397 77344 170812 77346
rect 170397 77288 170402 77344
rect 170458 77288 170812 77344
rect 170397 77286 170812 77288
rect 170397 77283 170463 77286
rect 170806 77284 170812 77286
rect 170876 77284 170882 77348
rect 143809 77210 143875 77213
rect 138430 77208 143875 77210
rect 138430 77152 143814 77208
rect 143870 77152 143875 77208
rect 138430 77150 143875 77152
rect 143809 77147 143875 77150
rect 147581 77210 147647 77213
rect 282913 77210 282979 77213
rect 147581 77208 282979 77210
rect 147581 77152 147586 77208
rect 147642 77152 282918 77208
rect 282974 77152 282979 77208
rect 147581 77150 282979 77152
rect 147581 77147 147647 77150
rect 282913 77147 282979 77150
rect 136214 77012 136220 77076
rect 136284 77074 136290 77076
rect 141969 77074 142035 77077
rect 136284 77072 142035 77074
rect 136284 77016 141974 77072
rect 142030 77016 142035 77072
rect 136284 77014 142035 77016
rect 136284 77012 136290 77014
rect 141969 77011 142035 77014
rect 153142 77012 153148 77076
rect 153212 77074 153218 77076
rect 354673 77074 354739 77077
rect 153212 77072 354739 77074
rect 153212 77016 354678 77072
rect 354734 77016 354739 77072
rect 153212 77014 354739 77016
rect 153212 77012 153218 77014
rect 354673 77011 354739 77014
rect 155861 76938 155927 76941
rect 389173 76938 389239 76941
rect 155861 76936 389239 76938
rect 155861 76880 155866 76936
rect 155922 76880 389178 76936
rect 389234 76880 389239 76936
rect 155861 76878 389239 76880
rect 155861 76875 155927 76878
rect 389173 76875 389239 76878
rect 111793 76802 111859 76805
rect 134333 76802 134399 76805
rect 111793 76800 134399 76802
rect 111793 76744 111798 76800
rect 111854 76744 134338 76800
rect 134394 76744 134399 76800
rect 111793 76742 134399 76744
rect 111793 76739 111859 76742
rect 134333 76739 134399 76742
rect 148358 76740 148364 76804
rect 148428 76802 148434 76804
rect 148685 76802 148751 76805
rect 148428 76800 148751 76802
rect 148428 76744 148690 76800
rect 148746 76744 148751 76800
rect 148428 76742 148751 76744
rect 148428 76740 148434 76742
rect 148685 76739 148751 76742
rect 161381 76802 161447 76805
rect 459553 76802 459619 76805
rect 161381 76800 459619 76802
rect 161381 76744 161386 76800
rect 161442 76744 459558 76800
rect 459614 76744 459619 76800
rect 161381 76742 459619 76744
rect 161381 76739 161447 76742
rect 459553 76739 459619 76742
rect 37273 76666 37339 76669
rect 128445 76666 128511 76669
rect 37273 76664 128511 76666
rect 37273 76608 37278 76664
rect 37334 76608 128450 76664
rect 128506 76608 128511 76664
rect 37273 76606 128511 76608
rect 37273 76603 37339 76606
rect 128445 76603 128511 76606
rect 143022 76604 143028 76668
rect 143092 76666 143098 76668
rect 143257 76666 143323 76669
rect 143092 76664 143323 76666
rect 143092 76608 143262 76664
rect 143318 76608 143323 76664
rect 143092 76606 143323 76608
rect 143092 76604 143098 76606
rect 143257 76603 143323 76606
rect 143809 76666 143875 76669
rect 144126 76666 144132 76668
rect 143809 76664 144132 76666
rect 143809 76608 143814 76664
rect 143870 76608 144132 76664
rect 143809 76606 144132 76608
rect 143809 76603 143875 76606
rect 144126 76604 144132 76606
rect 144196 76604 144202 76668
rect 148041 76666 148107 76669
rect 148174 76666 148180 76668
rect 148041 76664 148180 76666
rect 148041 76608 148046 76664
rect 148102 76608 148180 76664
rect 148041 76606 148180 76608
rect 148041 76603 148107 76606
rect 148174 76604 148180 76606
rect 148244 76604 148250 76668
rect 148777 76666 148843 76669
rect 148910 76666 148916 76668
rect 148777 76664 148916 76666
rect 148777 76608 148782 76664
rect 148838 76608 148916 76664
rect 148777 76606 148916 76608
rect 148777 76603 148843 76606
rect 148910 76604 148916 76606
rect 148980 76604 148986 76668
rect 157926 76604 157932 76668
rect 157996 76666 158002 76668
rect 158437 76666 158503 76669
rect 157996 76664 158503 76666
rect 157996 76608 158442 76664
rect 158498 76608 158503 76664
rect 157996 76606 158503 76608
rect 157996 76604 158002 76606
rect 158437 76603 158503 76606
rect 165153 76666 165219 76669
rect 505093 76666 505159 76669
rect 165153 76664 505159 76666
rect 165153 76608 165158 76664
rect 165214 76608 505098 76664
rect 505154 76608 505159 76664
rect 165153 76606 505159 76608
rect 165153 76603 165219 76606
rect 505093 76603 505159 76606
rect 20713 76530 20779 76533
rect 127157 76530 127223 76533
rect 20713 76528 127223 76530
rect 20713 76472 20718 76528
rect 20774 76472 127162 76528
rect 127218 76472 127223 76528
rect 20713 76470 127223 76472
rect 20713 76467 20779 76470
rect 127157 76467 127223 76470
rect 169661 76530 169727 76533
rect 565813 76530 565879 76533
rect 169661 76528 565879 76530
rect 169661 76472 169666 76528
rect 169722 76472 565818 76528
rect 565874 76472 565879 76528
rect 169661 76470 565879 76472
rect 169661 76467 169727 76470
rect 565813 76467 565879 76470
rect 141785 76394 141851 76397
rect 173157 76394 173223 76397
rect 141785 76392 173223 76394
rect 141785 76336 141790 76392
rect 141846 76336 173162 76392
rect 173218 76336 173223 76392
rect 141785 76334 173223 76336
rect 141785 76331 141851 76334
rect 173157 76331 173223 76334
rect 144862 76196 144868 76260
rect 144932 76258 144938 76260
rect 147305 76258 147371 76261
rect 144932 76256 147371 76258
rect 144932 76200 147310 76256
rect 147366 76200 147371 76256
rect 144932 76198 147371 76200
rect 144932 76196 144938 76198
rect 147305 76195 147371 76198
rect 162853 76258 162919 76261
rect 171726 76258 171732 76260
rect 162853 76256 171732 76258
rect 162853 76200 162858 76256
rect 162914 76200 171732 76256
rect 162853 76198 171732 76200
rect 162853 76195 162919 76198
rect 171726 76196 171732 76198
rect 171796 76196 171802 76260
rect 166758 76060 166764 76124
rect 166828 76122 166834 76124
rect 166901 76122 166967 76125
rect 166828 76120 166967 76122
rect 166828 76064 166906 76120
rect 166962 76064 166967 76120
rect 166828 76062 166967 76064
rect 166828 76060 166834 76062
rect 166901 76059 166967 76062
rect 139393 75986 139459 75989
rect 139526 75986 139532 75988
rect 139393 75984 139532 75986
rect 139393 75928 139398 75984
rect 139454 75928 139532 75984
rect 139393 75926 139532 75928
rect 139393 75923 139459 75926
rect 139526 75924 139532 75926
rect 139596 75924 139602 75988
rect 144913 75986 144979 75989
rect 145046 75986 145052 75988
rect 144913 75984 145052 75986
rect 144913 75928 144918 75984
rect 144974 75928 145052 75984
rect 144913 75926 145052 75928
rect 144913 75923 144979 75926
rect 145046 75924 145052 75926
rect 145116 75924 145122 75988
rect 146886 75924 146892 75988
rect 146956 75986 146962 75988
rect 147489 75986 147555 75989
rect 146956 75984 147555 75986
rect 146956 75928 147494 75984
rect 147550 75928 147555 75984
rect 146956 75926 147555 75928
rect 146956 75924 146962 75926
rect 147489 75923 147555 75926
rect 159030 75924 159036 75988
rect 159100 75986 159106 75988
rect 160185 75986 160251 75989
rect 159100 75984 160251 75986
rect 159100 75928 160190 75984
rect 160246 75928 160251 75984
rect 159100 75926 160251 75928
rect 159100 75924 159106 75926
rect 160185 75923 160251 75926
rect 160369 75986 160435 75989
rect 160502 75986 160508 75988
rect 160369 75984 160508 75986
rect 160369 75928 160374 75984
rect 160430 75928 160508 75984
rect 160369 75926 160508 75928
rect 160369 75923 160435 75926
rect 160502 75924 160508 75926
rect 160572 75924 160578 75988
rect 162342 75924 162348 75988
rect 162412 75986 162418 75988
rect 162761 75986 162827 75989
rect 165337 75988 165403 75989
rect 165286 75986 165292 75988
rect 162412 75984 162827 75986
rect 162412 75928 162766 75984
rect 162822 75928 162827 75984
rect 162412 75926 162827 75928
rect 165246 75926 165292 75986
rect 165356 75984 165403 75988
rect 165981 75988 166047 75989
rect 165981 75986 166028 75988
rect 165398 75928 165403 75984
rect 162412 75924 162418 75926
rect 162761 75923 162827 75926
rect 165286 75924 165292 75926
rect 165356 75924 165403 75928
rect 165936 75984 166028 75986
rect 165936 75928 165986 75984
rect 165936 75926 166028 75928
rect 165337 75923 165403 75924
rect 165981 75924 166028 75926
rect 166092 75924 166098 75988
rect 166206 75924 166212 75988
rect 166276 75986 166282 75988
rect 166533 75986 166599 75989
rect 166276 75984 166599 75986
rect 166276 75928 166538 75984
rect 166594 75928 166599 75984
rect 166276 75926 166599 75928
rect 166276 75924 166282 75926
rect 165981 75923 166047 75924
rect 166533 75923 166599 75926
rect 167310 75924 167316 75988
rect 167380 75986 167386 75988
rect 168005 75986 168071 75989
rect 167380 75984 168071 75986
rect 167380 75928 168010 75984
rect 168066 75928 168071 75984
rect 167380 75926 168071 75928
rect 167380 75924 167386 75926
rect 168005 75923 168071 75926
rect 140078 75788 140084 75852
rect 140148 75850 140154 75852
rect 140589 75850 140655 75853
rect 140148 75848 140655 75850
rect 140148 75792 140594 75848
rect 140650 75792 140655 75848
rect 140148 75790 140655 75792
rect 140148 75788 140154 75790
rect 140589 75787 140655 75790
rect 145414 75788 145420 75852
rect 145484 75850 145490 75852
rect 146017 75850 146083 75853
rect 145484 75848 146083 75850
rect 145484 75792 146022 75848
rect 146078 75792 146083 75848
rect 145484 75790 146083 75792
rect 145484 75788 145490 75790
rect 146017 75787 146083 75790
rect 160645 75850 160711 75853
rect 160870 75850 160876 75852
rect 160645 75848 160876 75850
rect 160645 75792 160650 75848
rect 160706 75792 160876 75848
rect 160645 75790 160876 75792
rect 160645 75787 160711 75790
rect 160870 75788 160876 75790
rect 160940 75788 160946 75852
rect 161790 75788 161796 75852
rect 161860 75850 161866 75852
rect 162025 75850 162091 75853
rect 161860 75848 162091 75850
rect 161860 75792 162030 75848
rect 162086 75792 162091 75848
rect 161860 75790 162091 75792
rect 161860 75788 161866 75790
rect 162025 75787 162091 75790
rect 162393 75850 162459 75853
rect 180057 75850 180123 75853
rect 162393 75848 180123 75850
rect 162393 75792 162398 75848
rect 162454 75792 180062 75848
rect 180118 75792 180123 75848
rect 162393 75790 180123 75792
rect 162393 75787 162459 75790
rect 180057 75787 180123 75790
rect 139158 75652 139164 75716
rect 139228 75714 139234 75716
rect 173893 75714 173959 75717
rect 139228 75712 173959 75714
rect 139228 75656 173898 75712
rect 173954 75656 173959 75712
rect 139228 75654 173959 75656
rect 139228 75652 139234 75654
rect 173893 75651 173959 75654
rect 140681 75578 140747 75581
rect 194593 75578 194659 75581
rect 140681 75576 194659 75578
rect 140681 75520 140686 75576
rect 140742 75520 194598 75576
rect 194654 75520 194659 75576
rect 140681 75518 194659 75520
rect 140681 75515 140747 75518
rect 194593 75515 194659 75518
rect 157149 75442 157215 75445
rect 402973 75442 403039 75445
rect 157149 75440 403039 75442
rect 157149 75384 157154 75440
rect 157210 75384 402978 75440
rect 403034 75384 403039 75440
rect 157149 75382 403039 75384
rect 157149 75379 157215 75382
rect 402973 75379 403039 75382
rect 2773 75306 2839 75309
rect 123661 75306 123727 75309
rect 2773 75304 123727 75306
rect 2773 75248 2778 75304
rect 2834 75248 123666 75304
rect 123722 75248 123727 75304
rect 2773 75246 123727 75248
rect 2773 75243 2839 75246
rect 123661 75243 123727 75246
rect 156229 75306 156295 75309
rect 164141 75306 164207 75309
rect 496813 75306 496879 75309
rect 156229 75304 156338 75306
rect 156229 75248 156234 75304
rect 156290 75248 156338 75304
rect 156229 75243 156338 75248
rect 164141 75304 496879 75306
rect 164141 75248 164146 75304
rect 164202 75248 496818 75304
rect 496874 75248 496879 75304
rect 164141 75246 496879 75248
rect 164141 75243 164207 75246
rect 496813 75243 496879 75246
rect 1393 75170 1459 75173
rect 125593 75170 125659 75173
rect 1393 75168 125659 75170
rect 1393 75112 1398 75168
rect 1454 75112 125598 75168
rect 125654 75112 125659 75168
rect 1393 75110 125659 75112
rect 156278 75170 156338 75243
rect 156689 75170 156755 75173
rect 156278 75168 156755 75170
rect 156278 75112 156694 75168
rect 156750 75112 156755 75168
rect 156278 75110 156755 75112
rect 1393 75107 1459 75110
rect 125593 75107 125659 75110
rect 156689 75107 156755 75110
rect 168281 75170 168347 75173
rect 549253 75170 549319 75173
rect 168281 75168 549319 75170
rect 168281 75112 168286 75168
rect 168342 75112 549258 75168
rect 549314 75112 549319 75168
rect 168281 75110 549319 75112
rect 168281 75107 168347 75110
rect 549253 75107 549319 75110
rect 161422 74972 161428 75036
rect 161492 75034 161498 75036
rect 171910 75034 171916 75036
rect 161492 74974 171916 75034
rect 161492 74972 161498 74974
rect 171910 74972 171916 74974
rect 171980 74972 171986 75036
rect 130377 74490 130443 74493
rect 135294 74490 135300 74492
rect 130377 74488 135300 74490
rect 130377 74432 130382 74488
rect 130438 74432 135300 74488
rect 130377 74430 135300 74432
rect 130377 74427 130443 74430
rect 135294 74428 135300 74430
rect 135364 74428 135370 74492
rect 158110 74428 158116 74492
rect 158180 74490 158186 74492
rect 158345 74490 158411 74493
rect 158180 74488 158411 74490
rect 158180 74432 158350 74488
rect 158406 74432 158411 74488
rect 158180 74430 158411 74432
rect 158180 74428 158186 74430
rect 158345 74427 158411 74430
rect 71773 74218 71839 74221
rect 131062 74218 131068 74220
rect 71773 74216 131068 74218
rect 71773 74160 71778 74216
rect 71834 74160 131068 74216
rect 71773 74158 131068 74160
rect 71773 74155 71839 74158
rect 131062 74156 131068 74158
rect 131132 74156 131138 74220
rect 145230 74156 145236 74220
rect 145300 74218 145306 74220
rect 146201 74218 146267 74221
rect 145300 74216 146267 74218
rect 145300 74160 146206 74216
rect 146262 74160 146267 74216
rect 145300 74158 146267 74160
rect 145300 74156 145306 74158
rect 146201 74155 146267 74158
rect 57973 74082 58039 74085
rect 130326 74082 130332 74084
rect 57973 74080 130332 74082
rect 57973 74024 57978 74080
rect 58034 74024 130332 74080
rect 57973 74022 130332 74024
rect 57973 74019 58039 74022
rect 130326 74020 130332 74022
rect 130396 74020 130402 74084
rect 143441 74082 143507 74085
rect 230473 74082 230539 74085
rect 143441 74080 230539 74082
rect 143441 74024 143446 74080
rect 143502 74024 230478 74080
rect 230534 74024 230539 74080
rect 143441 74022 230539 74024
rect 143441 74019 143507 74022
rect 230473 74019 230539 74022
rect 53833 73946 53899 73949
rect 130142 73946 130148 73948
rect 53833 73944 130148 73946
rect 53833 73888 53838 73944
rect 53894 73888 130148 73944
rect 53833 73886 130148 73888
rect 53833 73883 53899 73886
rect 130142 73884 130148 73886
rect 130212 73884 130218 73948
rect 144637 73946 144703 73949
rect 244273 73946 244339 73949
rect 144637 73944 244339 73946
rect 144637 73888 144642 73944
rect 144698 73888 244278 73944
rect 244334 73888 244339 73944
rect 144637 73886 244339 73888
rect 144637 73883 144703 73886
rect 244273 73883 244339 73886
rect 35893 73810 35959 73813
rect 128854 73810 128860 73812
rect 35893 73808 128860 73810
rect 35893 73752 35898 73808
rect 35954 73752 128860 73808
rect 35893 73750 128860 73752
rect 35893 73747 35959 73750
rect 128854 73748 128860 73750
rect 128924 73748 128930 73812
rect 170438 73748 170444 73812
rect 170508 73810 170514 73812
rect 578233 73810 578299 73813
rect 170508 73808 578299 73810
rect 170508 73752 578238 73808
rect 578294 73752 578299 73808
rect 170508 73750 578299 73752
rect 170508 73748 170514 73750
rect 578233 73747 578299 73750
rect 166206 73204 166212 73268
rect 166276 73266 166282 73268
rect 166717 73266 166783 73269
rect 166276 73264 166783 73266
rect 166276 73208 166722 73264
rect 166778 73208 166783 73264
rect 166276 73206 166783 73208
rect 166276 73204 166282 73206
rect 166717 73203 166783 73206
rect 140262 73068 140268 73132
rect 140332 73130 140338 73132
rect 140497 73130 140563 73133
rect 140332 73128 140563 73130
rect 140332 73072 140502 73128
rect 140558 73072 140563 73128
rect 140332 73070 140563 73072
rect 140332 73068 140338 73070
rect 140497 73067 140563 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 148910 72524 148916 72588
rect 148980 72586 148986 72588
rect 298093 72586 298159 72589
rect 148980 72584 298159 72586
rect 148980 72528 298098 72584
rect 298154 72528 298159 72584
rect 148980 72526 298159 72528
rect 148980 72524 148986 72526
rect 298093 72523 298159 72526
rect 172278 72388 172284 72452
rect 172348 72450 172354 72452
rect 500953 72450 501019 72453
rect 172348 72448 501019 72450
rect 172348 72392 500958 72448
rect 501014 72392 501019 72448
rect 172348 72390 501019 72392
rect 172348 72388 172354 72390
rect 500953 72387 501019 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 138790 69532 138796 69596
rect 138860 69594 138866 69596
rect 173249 69594 173315 69597
rect 138860 69592 173315 69594
rect 138860 69536 173254 69592
rect 173310 69536 173315 69592
rect 138860 69534 173315 69536
rect 138860 69532 138866 69534
rect 173249 69531 173315 69534
rect 152590 68172 152596 68236
rect 152660 68234 152666 68236
rect 353293 68234 353359 68237
rect 152660 68232 353359 68234
rect 152660 68176 353298 68232
rect 353354 68176 353359 68232
rect 152660 68174 353359 68176
rect 152660 68172 152666 68174
rect 353293 68171 353359 68174
rect 166206 66812 166212 66876
rect 166276 66874 166282 66876
rect 529933 66874 529999 66877
rect 166276 66872 529999 66874
rect 166276 66816 529938 66872
rect 529994 66816 529999 66872
rect 166276 66814 529999 66816
rect 166276 66812 166282 66814
rect 529933 66811 529999 66814
rect 140262 65452 140268 65516
rect 140332 65514 140338 65516
rect 193213 65514 193279 65517
rect 140332 65512 193279 65514
rect 140332 65456 193218 65512
rect 193274 65456 193279 65512
rect 140332 65454 193279 65456
rect 140332 65452 140338 65454
rect 193213 65451 193279 65454
rect 138974 62732 138980 62796
rect 139044 62794 139050 62796
rect 176653 62794 176719 62797
rect 139044 62792 176719 62794
rect 139044 62736 176658 62792
rect 176714 62736 176719 62792
rect 139044 62734 176719 62736
rect 139044 62732 139050 62734
rect 176653 62731 176719 62734
rect 138606 61372 138612 61436
rect 138676 61434 138682 61436
rect 172513 61434 172579 61437
rect 138676 61432 172579 61434
rect 138676 61376 172518 61432
rect 172574 61376 172579 61432
rect 138676 61374 172579 61376
rect 138676 61372 138682 61374
rect 172513 61371 172579 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 153878 58516 153884 58580
rect 153948 58578 153954 58580
rect 372613 58578 372679 58581
rect 153948 58576 372679 58578
rect 153948 58520 372618 58576
rect 372674 58520 372679 58576
rect 153948 58518 372679 58520
rect 153948 58516 153954 58518
rect 372613 58515 372679 58518
rect 165102 55796 165108 55860
rect 165172 55858 165178 55860
rect 511993 55858 512059 55861
rect 165172 55856 512059 55858
rect 165172 55800 511998 55856
rect 512054 55800 512059 55856
rect 165172 55798 512059 55800
rect 165172 55796 165178 55798
rect 511993 55795 512059 55798
rect 152774 51716 152780 51780
rect 152844 51778 152850 51780
rect 351913 51778 351979 51781
rect 152844 51776 351979 51778
rect 152844 51720 351918 51776
rect 351974 51720 351979 51776
rect 152844 51718 351979 51720
rect 152844 51716 152850 51718
rect 351913 51715 351979 51718
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 91093 44842 91159 44845
rect 133270 44842 133276 44844
rect 91093 44840 133276 44842
rect 91093 44784 91098 44840
rect 91154 44784 133276 44840
rect 91093 44782 133276 44784
rect 91093 44779 91159 44782
rect 133270 44780 133276 44782
rect 133340 44780 133346 44844
rect 172094 42060 172100 42124
rect 172164 42122 172170 42124
rect 550633 42122 550699 42125
rect 172164 42120 550699 42122
rect 172164 42064 550638 42120
rect 550694 42064 550699 42120
rect 172164 42062 550699 42064
rect 172164 42060 172170 42062
rect 550633 42059 550699 42062
rect 149462 35260 149468 35324
rect 149532 35322 149538 35324
rect 316033 35322 316099 35325
rect 149532 35320 316099 35322
rect 149532 35264 316038 35320
rect 316094 35264 316099 35320
rect 149532 35262 316099 35264
rect 149532 35260 149538 35262
rect 316033 35259 316099 35262
rect 163446 35124 163452 35188
rect 163516 35186 163522 35188
rect 473997 35186 474063 35189
rect 163516 35184 474063 35186
rect 163516 35128 474002 35184
rect 474058 35128 474063 35184
rect 163516 35126 474063 35128
rect 163516 35124 163522 35126
rect 473997 35123 474063 35126
rect 140998 34036 141004 34100
rect 141068 34098 141074 34100
rect 212533 34098 212599 34101
rect 141068 34096 212599 34098
rect 141068 34040 212538 34096
rect 212594 34040 212599 34096
rect 141068 34038 212599 34040
rect 141068 34036 141074 34038
rect 212533 34035 212599 34038
rect 143022 33900 143028 33964
rect 143092 33962 143098 33964
rect 226425 33962 226491 33965
rect 143092 33960 226491 33962
rect 143092 33904 226430 33960
rect 226486 33904 226491 33960
rect 143092 33902 226491 33904
rect 143092 33900 143098 33902
rect 226425 33899 226491 33902
rect 145230 33764 145236 33828
rect 145300 33826 145306 33828
rect 266353 33826 266419 33829
rect 145300 33824 266419 33826
rect 145300 33768 266358 33824
rect 266414 33768 266419 33824
rect 145300 33766 266419 33768
rect 145300 33764 145306 33766
rect 266353 33763 266419 33766
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 151302 31044 151308 31108
rect 151372 31106 151378 31108
rect 336733 31106 336799 31109
rect 151372 31104 336799 31106
rect 151372 31048 336738 31104
rect 336794 31048 336799 31104
rect 151372 31046 336799 31048
rect 151372 31044 151378 31046
rect 336733 31043 336799 31046
rect 169518 30908 169524 30972
rect 169588 30970 169594 30972
rect 567193 30970 567259 30973
rect 169588 30968 567259 30970
rect 169588 30912 567198 30968
rect 567254 30912 567259 30968
rect 169588 30910 567259 30912
rect 169588 30908 169594 30910
rect 567193 30907 567259 30910
rect 157926 29548 157932 29612
rect 157996 29610 158002 29612
rect 422293 29610 422359 29613
rect 157996 29608 422359 29610
rect 157996 29552 422298 29608
rect 422354 29552 422359 29608
rect 157996 29550 422359 29552
rect 157996 29548 158002 29550
rect 422293 29547 422359 29550
rect 151486 28324 151492 28388
rect 151556 28386 151562 28388
rect 335353 28386 335419 28389
rect 151556 28384 335419 28386
rect 151556 28328 335358 28384
rect 335414 28328 335419 28384
rect 151556 28326 335419 28328
rect 151556 28324 151562 28326
rect 335353 28323 335419 28326
rect 166390 28188 166396 28252
rect 166460 28250 166466 28252
rect 531313 28250 531379 28253
rect 166460 28248 531379 28250
rect 166460 28192 531318 28248
rect 531374 28192 531379 28248
rect 166460 28190 531379 28192
rect 166460 28188 166466 28190
rect 531313 28187 531379 28190
rect 144310 26964 144316 27028
rect 144380 27026 144386 27028
rect 242893 27026 242959 27029
rect 144380 27024 242959 27026
rect 144380 26968 242898 27024
rect 242954 26968 242959 27024
rect 144380 26966 242959 26968
rect 144380 26964 144386 26966
rect 242893 26963 242959 26966
rect 149646 26828 149652 26892
rect 149716 26890 149722 26892
rect 317413 26890 317479 26893
rect 149716 26888 317479 26890
rect 149716 26832 317418 26888
rect 317474 26832 317479 26888
rect 149716 26830 317479 26832
rect 149716 26828 149722 26830
rect 317413 26827 317479 26830
rect 162342 22748 162348 22812
rect 162412 22810 162418 22812
rect 477493 22810 477559 22813
rect 162412 22808 477559 22810
rect 162412 22752 477498 22808
rect 477554 22752 477559 22808
rect 162412 22750 477559 22752
rect 162412 22748 162418 22750
rect 477493 22747 477559 22750
rect 170622 22612 170628 22676
rect 170692 22674 170698 22676
rect 582373 22674 582439 22677
rect 170692 22672 582439 22674
rect 170692 22616 582378 22672
rect 582434 22616 582439 22672
rect 170692 22614 582439 22616
rect 170692 22612 170698 22614
rect 582373 22611 582439 22614
rect 159030 21252 159036 21316
rect 159100 21314 159106 21316
rect 442993 21314 443059 21317
rect 159100 21312 443059 21314
rect 159100 21256 442998 21312
rect 443054 21256 443059 21312
rect 159100 21254 443059 21256
rect 159100 21252 159106 21254
rect 442993 21251 443059 21254
rect 144494 20436 144500 20500
rect 144564 20498 144570 20500
rect 248413 20498 248479 20501
rect 144564 20496 248479 20498
rect 144564 20440 248418 20496
rect 248474 20440 248479 20496
rect 144564 20438 248479 20440
rect 144564 20436 144570 20438
rect 248413 20435 248479 20438
rect 156822 20300 156828 20364
rect 156892 20362 156898 20364
rect 407113 20362 407179 20365
rect 156892 20360 407179 20362
rect 156892 20304 407118 20360
rect 407174 20304 407179 20360
rect 156892 20302 407179 20304
rect 156892 20300 156898 20302
rect 407113 20299 407179 20302
rect 161054 20164 161060 20228
rect 161124 20226 161130 20228
rect 456793 20226 456859 20229
rect 161124 20224 456859 20226
rect 161124 20168 456798 20224
rect 456854 20168 456859 20224
rect 161124 20166 456859 20168
rect 161124 20164 161130 20166
rect 456793 20163 456859 20166
rect 160686 20028 160692 20092
rect 160756 20090 160762 20092
rect 458173 20090 458239 20093
rect 160756 20088 458239 20090
rect 160756 20032 458178 20088
rect 458234 20032 458239 20088
rect 160756 20030 458239 20032
rect 160756 20028 160762 20030
rect 458173 20027 458239 20030
rect 162526 19892 162532 19956
rect 162596 19954 162602 19956
rect 476113 19954 476179 19957
rect 162596 19952 476179 19954
rect 162596 19896 476118 19952
rect 476174 19896 476179 19952
rect 162596 19894 476179 19896
rect 162596 19892 162602 19894
rect 476113 19891 476179 19894
rect 579613 19818 579679 19821
rect 583520 19818 584960 19908
rect 579613 19816 584960 19818
rect 579613 19760 579618 19816
rect 579674 19760 584960 19816
rect 579613 19758 584960 19760
rect 579613 19755 579679 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3325 19410 3391 19413
rect -960 19408 3391 19410
rect -960 19352 3330 19408
rect 3386 19352 3391 19408
rect -960 19350 3391 19352
rect -960 19260 480 19350
rect 3325 19347 3391 19350
rect 166574 18668 166580 18732
rect 166644 18730 166650 18732
rect 531405 18730 531471 18733
rect 166644 18728 531471 18730
rect 166644 18672 531410 18728
rect 531466 18672 531471 18728
rect 166644 18670 531471 18672
rect 166644 18668 166650 18670
rect 531405 18667 531471 18670
rect 167678 18532 167684 18596
rect 167748 18594 167754 18596
rect 546493 18594 546559 18597
rect 167748 18592 546559 18594
rect 167748 18536 546498 18592
rect 546554 18536 546559 18592
rect 167748 18534 546559 18536
rect 167748 18532 167754 18534
rect 546493 18531 546559 18534
rect 134926 17852 134932 17916
rect 134996 17914 135002 17916
rect 251173 17914 251239 17917
rect 134996 17912 251239 17914
rect 134996 17856 251178 17912
rect 251234 17856 251239 17912
rect 134996 17854 251239 17856
rect 134996 17852 135002 17854
rect 251173 17851 251239 17854
rect 147070 17716 147076 17780
rect 147140 17778 147146 17780
rect 280153 17778 280219 17781
rect 147140 17776 280219 17778
rect 147140 17720 280158 17776
rect 280214 17720 280219 17776
rect 147140 17718 280219 17720
rect 147140 17716 147146 17718
rect 280153 17715 280219 17718
rect 136030 17580 136036 17644
rect 136100 17642 136106 17644
rect 284385 17642 284451 17645
rect 136100 17640 284451 17642
rect 136100 17584 284390 17640
rect 284446 17584 284451 17640
rect 136100 17582 284451 17584
rect 136100 17580 136106 17582
rect 284385 17579 284451 17582
rect 148542 17444 148548 17508
rect 148612 17506 148618 17508
rect 300853 17506 300919 17509
rect 148612 17504 300919 17506
rect 148612 17448 300858 17504
rect 300914 17448 300919 17504
rect 148612 17446 300919 17448
rect 148612 17444 148618 17446
rect 300853 17443 300919 17446
rect 157006 17308 157012 17372
rect 157076 17370 157082 17372
rect 405733 17370 405799 17373
rect 157076 17368 405799 17370
rect 157076 17312 405738 17368
rect 405794 17312 405799 17368
rect 157076 17310 405799 17312
rect 157076 17308 157082 17310
rect 405733 17307 405799 17310
rect 158110 17172 158116 17236
rect 158180 17234 158186 17236
rect 423673 17234 423739 17237
rect 158180 17232 423739 17234
rect 158180 17176 423678 17232
rect 423734 17176 423739 17232
rect 158180 17174 423739 17176
rect 158180 17172 158186 17174
rect 423673 17171 423739 17174
rect 140446 17036 140452 17100
rect 140516 17098 140522 17100
rect 191833 17098 191899 17101
rect 140516 17096 191899 17098
rect 140516 17040 191838 17096
rect 191894 17040 191899 17096
rect 140516 17038 191899 17040
rect 140516 17036 140522 17038
rect 191833 17035 191899 17038
rect 154062 16084 154068 16148
rect 154132 16146 154138 16148
rect 365713 16146 365779 16149
rect 154132 16144 365779 16146
rect 154132 16088 365718 16144
rect 365774 16088 365779 16144
rect 154132 16086 365779 16088
rect 154132 16084 154138 16086
rect 365713 16083 365779 16086
rect 155718 15948 155724 16012
rect 155788 16010 155794 16012
rect 387793 16010 387859 16013
rect 155788 16008 387859 16010
rect 155788 15952 387798 16008
rect 387854 15952 387859 16008
rect 155788 15950 387859 15952
rect 155788 15948 155794 15950
rect 387793 15947 387859 15950
rect 162710 15812 162716 15876
rect 162780 15874 162786 15876
rect 473353 15874 473419 15877
rect 162780 15872 473419 15874
rect 162780 15816 473358 15872
rect 473414 15816 473419 15872
rect 162780 15814 473419 15816
rect 162780 15812 162786 15814
rect 473353 15811 473419 15814
rect 145414 14860 145420 14924
rect 145484 14922 145490 14924
rect 264973 14922 265039 14925
rect 145484 14920 265039 14922
rect 145484 14864 264978 14920
rect 265034 14864 265039 14920
rect 145484 14862 265039 14864
rect 145484 14860 145490 14862
rect 264973 14859 265039 14862
rect 147254 14724 147260 14788
rect 147324 14786 147330 14788
rect 279049 14786 279115 14789
rect 147324 14784 279115 14786
rect 147324 14728 279054 14784
rect 279110 14728 279115 14784
rect 147324 14726 279115 14728
rect 147324 14724 147330 14726
rect 279049 14723 279115 14726
rect 154246 14588 154252 14652
rect 154316 14650 154322 14652
rect 370129 14650 370195 14653
rect 154316 14648 370195 14650
rect 154316 14592 370134 14648
rect 370190 14592 370195 14648
rect 154316 14590 370195 14592
rect 154316 14588 154322 14590
rect 370129 14587 370195 14590
rect 165286 14452 165292 14516
rect 165356 14514 165362 14516
rect 511257 14514 511323 14517
rect 165356 14512 511323 14514
rect 165356 14456 511262 14512
rect 511318 14456 511323 14512
rect 165356 14454 511323 14456
rect 165356 14452 165362 14454
rect 511257 14451 511323 14454
rect 143206 13228 143212 13292
rect 143276 13290 143282 13292
rect 229369 13290 229435 13293
rect 143276 13288 229435 13290
rect 143276 13232 229374 13288
rect 229430 13232 229435 13288
rect 143276 13230 229435 13232
rect 143276 13228 143282 13230
rect 229369 13227 229435 13230
rect 154430 13092 154436 13156
rect 154500 13154 154506 13156
rect 371233 13154 371299 13157
rect 154500 13152 371299 13154
rect 154500 13096 371238 13152
rect 371294 13096 371299 13152
rect 154500 13094 371299 13096
rect 154500 13092 154506 13094
rect 371233 13091 371299 13094
rect 166758 12956 166764 13020
rect 166828 13018 166834 13020
rect 528553 13018 528619 13021
rect 166828 13016 528619 13018
rect 166828 12960 528558 13016
rect 528614 12960 528619 13016
rect 166828 12958 528619 12960
rect 166828 12956 166834 12958
rect 528553 12955 528619 12958
rect 151670 12004 151676 12068
rect 151740 12066 151746 12068
rect 334617 12066 334683 12069
rect 151740 12064 334683 12066
rect 151740 12008 334622 12064
rect 334678 12008 334683 12064
rect 151740 12006 334683 12008
rect 151740 12004 151746 12006
rect 334617 12003 334683 12006
rect 158294 11868 158300 11932
rect 158364 11930 158370 11932
rect 423765 11930 423831 11933
rect 158364 11928 423831 11930
rect 158364 11872 423770 11928
rect 423826 11872 423831 11928
rect 158364 11870 423831 11872
rect 158364 11868 158370 11870
rect 423765 11867 423831 11870
rect 165470 11732 165476 11796
rect 165540 11794 165546 11796
rect 513373 11794 513439 11797
rect 165540 11792 513439 11794
rect 165540 11736 513378 11792
rect 513434 11736 513439 11792
rect 165540 11734 513439 11736
rect 165540 11732 165546 11734
rect 513373 11731 513439 11734
rect 169753 11658 169819 11661
rect 574645 11658 574711 11661
rect 169753 11656 574711 11658
rect 169753 11600 169758 11656
rect 169814 11600 574650 11656
rect 574706 11600 574711 11656
rect 169753 11598 574711 11600
rect 169753 11595 169819 11598
rect 574645 11595 574711 11598
rect 110505 10570 110571 10573
rect 134006 10570 134012 10572
rect 110505 10568 134012 10570
rect 110505 10512 110510 10568
rect 110566 10512 134012 10568
rect 110505 10510 134012 10512
rect 110505 10507 110571 10510
rect 134006 10508 134012 10510
rect 134076 10508 134082 10572
rect 92473 10434 92539 10437
rect 133086 10434 133092 10436
rect 92473 10432 133092 10434
rect 92473 10376 92478 10432
rect 92534 10376 133092 10432
rect 92473 10374 133092 10376
rect 92473 10371 92539 10374
rect 133086 10372 133092 10374
rect 133156 10372 133162 10436
rect 74993 10298 75059 10301
rect 131246 10298 131252 10300
rect 74993 10296 131252 10298
rect 74993 10240 74998 10296
rect 75054 10240 131252 10296
rect 74993 10238 131252 10240
rect 74993 10235 75059 10238
rect 131246 10236 131252 10238
rect 131316 10236 131322 10300
rect 158478 10236 158484 10300
rect 158548 10298 158554 10300
rect 420913 10298 420979 10301
rect 158548 10296 420979 10298
rect 158548 10240 420918 10296
rect 420974 10240 420979 10296
rect 158548 10238 420979 10240
rect 158548 10236 158554 10238
rect 420913 10235 420979 10238
rect 146886 9556 146892 9620
rect 146956 9618 146962 9620
rect 281901 9618 281967 9621
rect 146956 9616 281967 9618
rect 146956 9560 281906 9616
rect 281962 9560 281967 9616
rect 146956 9558 281967 9560
rect 146956 9556 146962 9558
rect 281901 9555 281967 9558
rect 148726 9420 148732 9484
rect 148796 9482 148802 9484
rect 299657 9482 299723 9485
rect 148796 9480 299723 9482
rect 148796 9424 299662 9480
rect 299718 9424 299723 9480
rect 148796 9422 299723 9424
rect 148796 9420 148802 9422
rect 299657 9419 299723 9422
rect 149830 9284 149836 9348
rect 149900 9346 149906 9348
rect 315021 9346 315087 9349
rect 149900 9344 315087 9346
rect 149900 9288 315026 9344
rect 315082 9288 315087 9344
rect 149900 9286 315087 9288
rect 149900 9284 149906 9286
rect 315021 9283 315087 9286
rect 57237 9210 57303 9213
rect 129958 9210 129964 9212
rect 57237 9208 129964 9210
rect 57237 9152 57242 9208
rect 57298 9152 129964 9208
rect 57237 9150 129964 9152
rect 57237 9147 57303 9150
rect 129958 9148 129964 9150
rect 130028 9148 130034 9212
rect 150014 9148 150020 9212
rect 150084 9210 150090 9212
rect 317321 9210 317387 9213
rect 150084 9208 317387 9210
rect 150084 9152 317326 9208
rect 317382 9152 317387 9208
rect 150084 9150 317387 9152
rect 150084 9148 150090 9150
rect 317321 9147 317387 9150
rect 56041 9074 56107 9077
rect 129774 9074 129780 9076
rect 56041 9072 129780 9074
rect 56041 9016 56046 9072
rect 56102 9016 129780 9072
rect 56041 9014 129780 9016
rect 56041 9011 56107 9014
rect 129774 9012 129780 9014
rect 129844 9012 129850 9076
rect 152406 9012 152412 9076
rect 152476 9074 152482 9076
rect 351637 9074 351703 9077
rect 152476 9072 351703 9074
rect 152476 9016 351642 9072
rect 351698 9016 351703 9072
rect 152476 9014 351703 9016
rect 152476 9012 152482 9014
rect 351637 9011 351703 9014
rect 41873 8938 41939 8941
rect 128670 8938 128676 8940
rect 41873 8936 128676 8938
rect 41873 8880 41878 8936
rect 41934 8880 128676 8936
rect 41873 8878 128676 8880
rect 41873 8875 41939 8878
rect 128670 8876 128676 8878
rect 128740 8876 128746 8940
rect 156638 8876 156644 8940
rect 156708 8938 156714 8940
rect 407205 8938 407271 8941
rect 156708 8936 407271 8938
rect 156708 8880 407210 8936
rect 407266 8880 407271 8936
rect 156708 8878 407271 8880
rect 156708 8876 156714 8878
rect 407205 8875 407271 8878
rect 133638 8740 133644 8804
rect 133708 8802 133714 8804
rect 197905 8802 197971 8805
rect 133708 8800 197971 8802
rect 133708 8744 197910 8800
rect 197966 8744 197971 8800
rect 133708 8742 197971 8744
rect 133708 8740 133714 8742
rect 197905 8739 197971 8742
rect 109309 7714 109375 7717
rect 134190 7714 134196 7716
rect 109309 7712 134196 7714
rect 109309 7656 109314 7712
rect 109370 7656 134196 7712
rect 109309 7654 134196 7656
rect 109309 7651 109375 7654
rect 134190 7652 134196 7654
rect 134260 7652 134266 7716
rect 23013 7578 23079 7581
rect 127198 7578 127204 7580
rect 23013 7576 127204 7578
rect 23013 7520 23018 7576
rect 23074 7520 127204 7576
rect 23013 7518 127204 7520
rect 23013 7515 23079 7518
rect 127198 7516 127204 7518
rect 127268 7516 127274 7580
rect 142838 6836 142844 6900
rect 142908 6898 142914 6900
rect 228725 6898 228791 6901
rect 142908 6896 228791 6898
rect 142908 6840 228730 6896
rect 228786 6840 228791 6896
rect 142908 6838 228791 6840
rect 142908 6836 142914 6838
rect 228725 6835 228791 6838
rect 144678 6700 144684 6764
rect 144748 6762 144754 6764
rect 246389 6762 246455 6765
rect 144748 6760 246455 6762
rect 144748 6704 246394 6760
rect 246450 6704 246455 6760
rect 144748 6702 246455 6704
rect 144748 6700 144754 6702
rect 246389 6699 246455 6702
rect -960 6490 480 6580
rect 145598 6564 145604 6628
rect 145668 6626 145674 6628
rect 264145 6626 264211 6629
rect 145668 6624 264211 6626
rect 145668 6568 264150 6624
rect 264206 6568 264211 6624
rect 145668 6566 264211 6568
rect 145668 6564 145674 6566
rect 264145 6563 264211 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 148358 6428 148364 6492
rect 148428 6490 148434 6492
rect 300761 6490 300827 6493
rect 148428 6488 300827 6490
rect 148428 6432 300766 6488
rect 300822 6432 300827 6488
rect 583520 6476 584960 6566
rect 148428 6430 300827 6432
rect 148428 6428 148434 6430
rect 300761 6427 300827 6430
rect 73797 6354 73863 6357
rect 131430 6354 131436 6356
rect 73797 6352 131436 6354
rect 73797 6296 73802 6352
rect 73858 6296 131436 6352
rect 73797 6294 131436 6296
rect 73797 6291 73863 6294
rect 131430 6292 131436 6294
rect 131500 6292 131506 6356
rect 167862 6292 167868 6356
rect 167932 6354 167938 6356
rect 549069 6354 549135 6357
rect 167932 6352 549135 6354
rect 167932 6296 549074 6352
rect 549130 6296 549135 6352
rect 167932 6294 549135 6296
rect 167932 6292 167938 6294
rect 549069 6291 549135 6294
rect 40677 6218 40743 6221
rect 128670 6218 128676 6220
rect 40677 6216 128676 6218
rect 40677 6160 40682 6216
rect 40738 6160 128676 6216
rect 40677 6158 128676 6160
rect 40677 6155 40743 6158
rect 128670 6156 128676 6158
rect 128740 6156 128746 6220
rect 137686 6156 137692 6220
rect 137756 6218 137762 6220
rect 160093 6218 160159 6221
rect 137756 6216 160159 6218
rect 137756 6160 160098 6216
rect 160154 6160 160159 6216
rect 137756 6158 160159 6160
rect 137756 6156 137762 6158
rect 160093 6155 160159 6158
rect 170806 6156 170812 6220
rect 170876 6218 170882 6220
rect 576301 6218 576367 6221
rect 170876 6216 576367 6218
rect 170876 6160 576306 6216
rect 576362 6160 576367 6216
rect 170876 6158 576367 6160
rect 170876 6156 170882 6158
rect 576301 6155 576367 6158
rect 140078 6020 140084 6084
rect 140148 6082 140154 6084
rect 194409 6082 194475 6085
rect 140148 6080 194475 6082
rect 140148 6024 194414 6080
rect 194470 6024 194475 6080
rect 140148 6022 194475 6024
rect 140148 6020 140154 6022
rect 194409 6019 194475 6022
rect 163630 5068 163636 5132
rect 163700 5130 163706 5132
rect 494697 5130 494763 5133
rect 163700 5128 494763 5130
rect 163700 5072 494702 5128
rect 494758 5072 494763 5128
rect 163700 5070 494763 5072
rect 163700 5068 163706 5070
rect 494697 5067 494763 5070
rect 168046 4932 168052 4996
rect 168116 4994 168122 4996
rect 547873 4994 547939 4997
rect 168116 4992 547939 4994
rect 168116 4936 547878 4992
rect 547934 4936 547939 4992
rect 168116 4934 547939 4936
rect 168116 4932 168122 4934
rect 547873 4931 547939 4934
rect 4061 4858 4127 4861
rect 125910 4858 125916 4860
rect 4061 4856 125916 4858
rect 4061 4800 4066 4856
rect 4122 4800 125916 4856
rect 4061 4798 125916 4800
rect 4061 4795 4127 4798
rect 125910 4796 125916 4798
rect 125980 4796 125986 4860
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 158897 4858 158963 4861
rect 137940 4856 158963 4858
rect 137940 4800 158902 4856
rect 158958 4800 158963 4856
rect 137940 4798 158963 4800
rect 137940 4796 137946 4798
rect 158897 4795 158963 4798
rect 170990 4796 170996 4860
rect 171060 4858 171066 4860
rect 577405 4858 577471 4861
rect 171060 4856 577471 4858
rect 171060 4800 577410 4856
rect 577466 4800 577471 4856
rect 171060 4798 577471 4800
rect 171060 4796 171066 4798
rect 577405 4795 577471 4798
rect 136398 3980 136404 4044
rect 136468 4042 136474 4044
rect 142429 4042 142495 4045
rect 136468 4040 142495 4042
rect 136468 3984 142434 4040
rect 142490 3984 142495 4040
rect 136468 3982 142495 3984
rect 136468 3980 136474 3982
rect 142429 3979 142495 3982
rect 146845 4042 146911 4045
rect 210969 4042 211035 4045
rect 146845 4040 211035 4042
rect 146845 3984 146850 4040
rect 146906 3984 210974 4040
rect 211030 3984 211035 4040
rect 146845 3982 211035 3984
rect 146845 3979 146911 3982
rect 210969 3979 211035 3982
rect 142337 3906 142403 3909
rect 218145 3906 218211 3909
rect 142337 3904 218211 3906
rect 142337 3848 142342 3904
rect 142398 3848 218150 3904
rect 218206 3848 218211 3904
rect 142337 3846 218211 3848
rect 142337 3843 142403 3846
rect 218145 3843 218211 3846
rect 131982 3708 131988 3772
rect 132052 3770 132058 3772
rect 221549 3770 221615 3773
rect 132052 3768 221615 3770
rect 132052 3712 221554 3768
rect 221610 3712 221615 3768
rect 132052 3710 221615 3712
rect 132052 3708 132058 3710
rect 221549 3707 221615 3710
rect 136214 3572 136220 3636
rect 136284 3634 136290 3636
rect 146845 3634 146911 3637
rect 235809 3634 235875 3637
rect 136284 3632 146911 3634
rect 136284 3576 146850 3632
rect 146906 3576 146911 3632
rect 136284 3574 146911 3576
rect 136284 3572 136290 3574
rect 146845 3571 146911 3574
rect 151770 3632 235875 3634
rect 151770 3576 235814 3632
rect 235870 3576 235875 3632
rect 151770 3574 235875 3576
rect 144545 3498 144611 3501
rect 151770 3498 151830 3574
rect 235809 3571 235875 3574
rect 144545 3496 151830 3498
rect 144545 3440 144550 3496
rect 144606 3440 151830 3496
rect 144545 3438 151830 3440
rect 144545 3435 144611 3438
rect 171910 3436 171916 3500
rect 171980 3498 171986 3500
rect 461577 3498 461643 3501
rect 171980 3496 461643 3498
rect 171980 3440 461582 3496
rect 461638 3440 461643 3496
rect 171980 3438 461643 3440
rect 171980 3436 171986 3438
rect 461577 3435 461643 3438
rect 20621 3362 20687 3365
rect 127382 3362 127388 3364
rect 20621 3360 127388 3362
rect 20621 3304 20626 3360
rect 20682 3304 127388 3360
rect 20621 3302 127388 3304
rect 20621 3299 20687 3302
rect 127382 3300 127388 3302
rect 127452 3300 127458 3364
rect 171726 3300 171732 3364
rect 171796 3362 171802 3364
rect 472249 3362 472315 3365
rect 171796 3360 472315 3362
rect 171796 3304 472254 3360
rect 472310 3304 472315 3360
rect 171796 3302 472315 3304
rect 171796 3300 171802 3302
rect 472249 3299 472315 3302
rect 143073 3226 143139 3229
rect 214465 3226 214531 3229
rect 143073 3224 214531 3226
rect 143073 3168 143078 3224
rect 143134 3168 214470 3224
rect 214526 3168 214531 3224
rect 143073 3166 214531 3168
rect 143073 3163 143139 3166
rect 214465 3163 214531 3166
<< via3 >>
rect 144132 187580 144196 187644
rect 140820 186280 140884 186284
rect 140820 186224 140834 186280
rect 140834 186224 140884 186280
rect 140820 186220 140884 186224
rect 143028 182684 143092 182748
rect 141556 182548 141620 182612
rect 141004 182412 141068 182476
rect 142476 180916 142540 180980
rect 146156 180916 146220 180980
rect 143028 178876 143092 178940
rect 141004 178740 141068 178804
rect 140820 178604 140884 178668
rect 141556 178468 141620 178532
rect 165476 175536 165540 175540
rect 165476 175480 165490 175536
rect 165490 175480 165540 175536
rect 165476 175476 165540 175480
rect 146156 174524 146220 174588
rect 142476 172952 142540 172956
rect 142476 172896 142526 172952
rect 142526 172896 142540 172952
rect 142476 172892 142540 172896
rect 165476 172952 165540 172956
rect 165476 172896 165490 172952
rect 165490 172896 165540 172952
rect 165476 172892 165540 172896
rect 144132 156572 144196 156636
rect 182220 141340 182284 141404
rect 118556 139980 118620 140044
rect 182220 110604 182284 110668
rect 118556 96324 118620 96388
rect 171364 80548 171428 80612
rect 129780 80004 129844 80068
rect 126284 79868 126348 79932
rect 127388 79868 127452 79932
rect 127756 79906 127760 79932
rect 127760 79906 127816 79932
rect 127816 79906 127820 79932
rect 127756 79868 127820 79906
rect 127388 79732 127452 79796
rect 128492 79868 128556 79932
rect 129228 79928 129292 79932
rect 141004 80140 141068 80204
rect 144868 80140 144932 80204
rect 152412 80140 152476 80204
rect 129228 79872 129232 79928
rect 129232 79872 129288 79928
rect 129288 79872 129292 79928
rect 129228 79868 129292 79872
rect 130884 79868 130948 79932
rect 130332 79732 130396 79796
rect 128676 79656 128740 79660
rect 128676 79600 128726 79656
rect 128726 79600 128740 79656
rect 128676 79596 128740 79600
rect 131252 79596 131316 79660
rect 132172 79906 132176 79932
rect 132176 79906 132232 79932
rect 132232 79906 132236 79932
rect 132172 79868 132236 79906
rect 133460 79868 133524 79932
rect 133092 79596 133156 79660
rect 135300 79732 135364 79796
rect 138060 79928 138124 79932
rect 138060 79872 138064 79928
rect 138064 79872 138120 79928
rect 138120 79872 138124 79928
rect 138060 79868 138124 79872
rect 139164 79868 139228 79932
rect 137876 79792 137940 79796
rect 137876 79736 137926 79792
rect 137926 79736 137940 79792
rect 137876 79732 137940 79736
rect 138980 79732 139044 79796
rect 140636 79868 140700 79932
rect 143212 79868 143276 79932
rect 144132 79906 144136 79932
rect 144136 79906 144192 79932
rect 144192 79906 144196 79932
rect 144132 79868 144196 79906
rect 141372 79732 141436 79796
rect 138612 79596 138676 79660
rect 139532 79656 139596 79660
rect 139532 79600 139582 79656
rect 139582 79600 139596 79656
rect 139532 79596 139596 79600
rect 142844 79732 142908 79796
rect 144684 79906 144688 79932
rect 144688 79906 144744 79932
rect 144744 79906 144748 79932
rect 144684 79868 144748 79906
rect 144316 79732 144380 79796
rect 144500 79732 144564 79796
rect 145420 80004 145484 80068
rect 145052 79868 145116 79932
rect 145604 79732 145668 79796
rect 147076 79868 147140 79932
rect 145420 79596 145484 79660
rect 147260 79792 147324 79796
rect 147260 79736 147310 79792
rect 147310 79736 147324 79792
rect 147260 79732 147324 79736
rect 163452 80140 163516 80204
rect 172284 80276 172348 80340
rect 148180 79868 148244 79932
rect 148732 79868 148796 79932
rect 148548 79732 148612 79796
rect 149652 79868 149716 79932
rect 150572 79868 150636 79932
rect 150020 79732 150084 79796
rect 151860 79928 151924 79932
rect 151860 79872 151864 79928
rect 151864 79872 151920 79928
rect 151920 79872 151924 79928
rect 151860 79868 151924 79872
rect 153148 79906 153152 79932
rect 153152 79906 153208 79932
rect 153208 79906 153212 79932
rect 153148 79868 153212 79906
rect 153884 79868 153948 79932
rect 155724 79928 155788 79932
rect 155724 79872 155728 79928
rect 155728 79872 155784 79928
rect 155784 79872 155788 79928
rect 155724 79868 155788 79872
rect 151492 79596 151556 79660
rect 152780 79732 152844 79796
rect 154068 79732 154132 79796
rect 154436 79792 154500 79796
rect 154436 79736 154486 79792
rect 154486 79736 154500 79792
rect 154436 79732 154500 79736
rect 154252 79596 154316 79660
rect 156828 79868 156892 79932
rect 156828 79596 156892 79660
rect 157932 79868 157996 79932
rect 158300 79928 158364 79932
rect 158300 79872 158304 79928
rect 158304 79872 158360 79928
rect 158360 79872 158364 79928
rect 158300 79868 158364 79872
rect 158300 79732 158364 79796
rect 157748 79596 157812 79660
rect 159956 79868 160020 79932
rect 160876 79928 160940 79932
rect 160876 79872 160880 79928
rect 160880 79872 160936 79928
rect 160936 79872 160940 79928
rect 160876 79868 160940 79872
rect 161060 79928 161124 79932
rect 161060 79872 161064 79928
rect 161064 79872 161120 79928
rect 161120 79872 161124 79928
rect 161060 79868 161124 79872
rect 161428 79906 161432 79932
rect 161432 79906 161488 79932
rect 161488 79906 161492 79932
rect 161428 79868 161492 79906
rect 161796 79868 161860 79932
rect 160508 79732 160572 79796
rect 162716 79732 162780 79796
rect 163084 79732 163148 79796
rect 165476 79928 165540 79932
rect 165476 79872 165480 79928
rect 165480 79872 165536 79928
rect 165536 79872 165540 79928
rect 165476 79868 165540 79872
rect 166028 79928 166092 79932
rect 166028 79872 166032 79928
rect 166032 79872 166088 79928
rect 166088 79872 166092 79928
rect 166028 79868 166092 79872
rect 166212 79928 166276 79932
rect 166212 79872 166216 79928
rect 166216 79872 166272 79928
rect 166272 79872 166276 79928
rect 166212 79868 166276 79872
rect 167316 79906 167320 79932
rect 167320 79906 167376 79932
rect 167376 79906 167380 79932
rect 167316 79868 167380 79906
rect 168052 79868 168116 79932
rect 166396 79732 166460 79796
rect 167684 79732 167748 79796
rect 172100 80140 172164 80204
rect 173020 80140 173084 80204
rect 169892 79928 169956 79932
rect 169892 79872 169896 79928
rect 169896 79872 169952 79928
rect 169952 79872 169956 79928
rect 160324 79596 160388 79660
rect 160692 79596 160756 79660
rect 162532 79596 162596 79660
rect 163268 79596 163332 79660
rect 163636 79596 163700 79660
rect 166580 79596 166644 79660
rect 169892 79868 169956 79872
rect 170812 79868 170876 79932
rect 171364 79906 171368 79932
rect 171368 79906 171424 79932
rect 171424 79906 171428 79932
rect 171364 79868 171428 79906
rect 171916 79868 171980 79932
rect 172652 79868 172716 79932
rect 173020 79928 173084 79932
rect 173020 79872 173024 79928
rect 173024 79872 173080 79928
rect 173080 79872 173084 79928
rect 173020 79868 173084 79872
rect 170628 79732 170692 79796
rect 172652 79732 172716 79796
rect 173388 79868 173452 79932
rect 173940 79928 174004 79932
rect 173940 79872 173944 79928
rect 173944 79872 174000 79928
rect 174000 79872 174004 79928
rect 173940 79868 174004 79872
rect 173572 79732 173636 79796
rect 169524 79596 169588 79660
rect 171916 79460 171980 79524
rect 172652 79460 172716 79524
rect 173388 79188 173452 79252
rect 128860 78780 128924 78844
rect 130148 78780 130212 78844
rect 136404 78780 136468 78844
rect 137692 78780 137756 78844
rect 140452 78780 140516 78844
rect 151308 78780 151372 78844
rect 159956 78780 160020 78844
rect 165108 78780 165172 78844
rect 172836 78780 172900 78844
rect 129228 78644 129292 78708
rect 129964 78704 130028 78708
rect 129964 78648 130014 78704
rect 130014 78648 130028 78704
rect 129964 78644 130028 78648
rect 131436 78644 131500 78708
rect 134012 78704 134076 78708
rect 134012 78648 134062 78704
rect 134062 78648 134076 78704
rect 134012 78644 134076 78648
rect 138060 78704 138124 78708
rect 138060 78648 138074 78704
rect 138074 78648 138124 78704
rect 138060 78644 138124 78648
rect 138796 78644 138860 78708
rect 151676 78644 151740 78708
rect 151860 78704 151924 78708
rect 151860 78648 151910 78704
rect 151910 78648 151924 78704
rect 151860 78644 151924 78648
rect 156644 78644 156708 78708
rect 160324 78644 160388 78708
rect 163268 78644 163332 78708
rect 173020 78644 173084 78708
rect 173204 78644 173268 78708
rect 173572 78508 173636 78572
rect 173940 78372 174004 78436
rect 133644 78236 133708 78300
rect 140636 78236 140700 78300
rect 132172 78100 132236 78164
rect 141372 78100 141436 78164
rect 149836 78100 149900 78164
rect 150572 78160 150636 78164
rect 150572 78104 150586 78160
rect 150586 78104 150636 78160
rect 150572 78100 150636 78104
rect 133276 77964 133340 78028
rect 134196 77964 134260 78028
rect 134932 77964 134996 78028
rect 125916 77828 125980 77892
rect 127572 77828 127636 77892
rect 133460 77828 133524 77892
rect 136036 77828 136100 77892
rect 138060 77828 138124 77892
rect 157932 77828 157996 77892
rect 126284 77692 126348 77756
rect 131988 77692 132052 77756
rect 168052 77420 168116 77484
rect 169892 77480 169956 77484
rect 169892 77424 169942 77480
rect 169942 77424 169956 77480
rect 169892 77420 169956 77424
rect 170444 77480 170508 77484
rect 170444 77424 170494 77480
rect 170494 77424 170508 77480
rect 170444 77420 170508 77424
rect 138060 77284 138124 77348
rect 149468 77284 149532 77348
rect 152596 77284 152660 77348
rect 157748 77344 157812 77348
rect 157748 77288 157798 77344
rect 157798 77288 157812 77344
rect 157748 77284 157812 77288
rect 163084 77284 163148 77348
rect 170812 77284 170876 77348
rect 136220 77012 136284 77076
rect 153148 77012 153212 77076
rect 148364 76740 148428 76804
rect 143028 76604 143092 76668
rect 144132 76604 144196 76668
rect 148180 76604 148244 76668
rect 148916 76604 148980 76668
rect 157932 76604 157996 76668
rect 144868 76196 144932 76260
rect 171732 76196 171796 76260
rect 166764 76060 166828 76124
rect 139532 75924 139596 75988
rect 145052 75924 145116 75988
rect 146892 75924 146956 75988
rect 159036 75924 159100 75988
rect 160508 75924 160572 75988
rect 162348 75924 162412 75988
rect 165292 75984 165356 75988
rect 165292 75928 165342 75984
rect 165342 75928 165356 75984
rect 165292 75924 165356 75928
rect 166028 75984 166092 75988
rect 166028 75928 166042 75984
rect 166042 75928 166092 75984
rect 166028 75924 166092 75928
rect 166212 75924 166276 75988
rect 167316 75924 167380 75988
rect 140084 75788 140148 75852
rect 145420 75788 145484 75852
rect 160876 75788 160940 75852
rect 161796 75788 161860 75852
rect 139164 75652 139228 75716
rect 161428 74972 161492 75036
rect 171916 74972 171980 75036
rect 135300 74428 135364 74492
rect 158116 74428 158180 74492
rect 131068 74156 131132 74220
rect 145236 74156 145300 74220
rect 130332 74020 130396 74084
rect 130148 73884 130212 73948
rect 128860 73748 128924 73812
rect 170444 73748 170508 73812
rect 166212 73204 166276 73268
rect 140268 73068 140332 73132
rect 148916 72524 148980 72588
rect 172284 72388 172348 72452
rect 138796 69532 138860 69596
rect 152596 68172 152660 68236
rect 166212 66812 166276 66876
rect 140268 65452 140332 65516
rect 138980 62732 139044 62796
rect 138612 61372 138676 61436
rect 153884 58516 153948 58580
rect 165108 55796 165172 55860
rect 152780 51716 152844 51780
rect 133276 44780 133340 44844
rect 172100 42060 172164 42124
rect 149468 35260 149532 35324
rect 163452 35124 163516 35188
rect 141004 34036 141068 34100
rect 143028 33900 143092 33964
rect 145236 33764 145300 33828
rect 151308 31044 151372 31108
rect 169524 30908 169588 30972
rect 157932 29548 157996 29612
rect 151492 28324 151556 28388
rect 166396 28188 166460 28252
rect 144316 26964 144380 27028
rect 149652 26828 149716 26892
rect 162348 22748 162412 22812
rect 170628 22612 170692 22676
rect 159036 21252 159100 21316
rect 144500 20436 144564 20500
rect 156828 20300 156892 20364
rect 161060 20164 161124 20228
rect 160692 20028 160756 20092
rect 162532 19892 162596 19956
rect 166580 18668 166644 18732
rect 167684 18532 167748 18596
rect 134932 17852 134996 17916
rect 147076 17716 147140 17780
rect 136036 17580 136100 17644
rect 148548 17444 148612 17508
rect 157012 17308 157076 17372
rect 158116 17172 158180 17236
rect 140452 17036 140516 17100
rect 154068 16084 154132 16148
rect 155724 15948 155788 16012
rect 162716 15812 162780 15876
rect 145420 14860 145484 14924
rect 147260 14724 147324 14788
rect 154252 14588 154316 14652
rect 165292 14452 165356 14516
rect 143212 13228 143276 13292
rect 154436 13092 154500 13156
rect 166764 12956 166828 13020
rect 151676 12004 151740 12068
rect 158300 11868 158364 11932
rect 165476 11732 165540 11796
rect 134012 10508 134076 10572
rect 133092 10372 133156 10436
rect 131252 10236 131316 10300
rect 158484 10236 158548 10300
rect 146892 9556 146956 9620
rect 148732 9420 148796 9484
rect 149836 9284 149900 9348
rect 129964 9148 130028 9212
rect 150020 9148 150084 9212
rect 129780 9012 129844 9076
rect 152412 9012 152476 9076
rect 128676 8876 128740 8940
rect 156644 8876 156708 8940
rect 133644 8740 133708 8804
rect 134196 7652 134260 7716
rect 127204 7516 127268 7580
rect 142844 6836 142908 6900
rect 144684 6700 144748 6764
rect 145604 6564 145668 6628
rect 148364 6428 148428 6492
rect 131436 6292 131500 6356
rect 167868 6292 167932 6356
rect 128676 6156 128740 6220
rect 137692 6156 137756 6220
rect 170812 6156 170876 6220
rect 140084 6020 140148 6084
rect 163636 5068 163700 5132
rect 168052 4932 168116 4996
rect 125916 4796 125980 4860
rect 137876 4796 137940 4860
rect 170996 4796 171060 4860
rect 136404 3980 136468 4044
rect 131988 3708 132052 3772
rect 136220 3572 136284 3636
rect 171916 3436 171980 3500
rect 127388 3300 127452 3364
rect 171732 3300 171796 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 144131 187644 144197 187645
rect 144131 187580 144132 187644
rect 144196 187580 144197 187644
rect 144131 187579 144197 187580
rect 140819 186284 140885 186285
rect 140819 186220 140820 186284
rect 140884 186220 140885 186284
rect 140819 186219 140885 186220
rect 140822 178669 140882 186219
rect 143027 182748 143093 182749
rect 143027 182684 143028 182748
rect 143092 182684 143093 182748
rect 143027 182683 143093 182684
rect 141555 182612 141621 182613
rect 141555 182548 141556 182612
rect 141620 182548 141621 182612
rect 141555 182547 141621 182548
rect 141003 182476 141069 182477
rect 141003 182412 141004 182476
rect 141068 182412 141069 182476
rect 141003 182411 141069 182412
rect 141006 178805 141066 182411
rect 141003 178804 141069 178805
rect 141003 178740 141004 178804
rect 141068 178740 141069 178804
rect 141003 178739 141069 178740
rect 140819 178668 140885 178669
rect 140819 178604 140820 178668
rect 140884 178604 140885 178668
rect 140819 178603 140885 178604
rect 141558 178533 141618 182547
rect 142475 180980 142541 180981
rect 142475 180916 142476 180980
rect 142540 180916 142541 180980
rect 142475 180915 142541 180916
rect 141555 178532 141621 178533
rect 141555 178468 141556 178532
rect 141620 178468 141621 178532
rect 141555 178467 141621 178468
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 142478 172957 142538 180915
rect 143030 178941 143090 182683
rect 143027 178940 143093 178941
rect 143027 178876 143028 178940
rect 143092 178876 143093 178940
rect 143027 178875 143093 178876
rect 142475 172956 142541 172957
rect 142475 172892 142476 172956
rect 142540 172892 142541 172956
rect 142475 172891 142541 172892
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 144134 156637 144194 187579
rect 146155 180980 146221 180981
rect 146155 180916 146156 180980
rect 146220 180916 146221 180980
rect 146155 180915 146221 180916
rect 146158 174589 146218 180915
rect 165475 175540 165541 175541
rect 165475 175476 165476 175540
rect 165540 175476 165541 175540
rect 165475 175475 165541 175476
rect 146155 174588 146221 174589
rect 146155 174524 146156 174588
rect 146220 174524 146221 174588
rect 146155 174523 146221 174524
rect 165478 172957 165538 175475
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 165475 172956 165541 172957
rect 165475 172892 165476 172956
rect 165540 172892 165541 172956
rect 165475 172891 165541 172892
rect 144131 156636 144197 156637
rect 144131 156572 144132 156636
rect 144196 156572 144197 156636
rect 144131 156571 144197 156572
rect 172794 142000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 182219 141404 182285 141405
rect 182219 141340 182220 141404
rect 182284 141340 182285 141404
rect 182219 141339 182285 141340
rect 118555 140044 118621 140045
rect 118555 139980 118556 140044
rect 118620 139980 118621 140044
rect 118555 139979 118621 139980
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 118558 96389 118618 139979
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 182222 110669 182282 141339
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 182219 110668 182285 110669
rect 182219 110604 182220 110668
rect 182284 110604 182285 110668
rect 182219 110603 182285 110604
rect 118555 96388 118621 96389
rect 118555 96324 118556 96388
rect 118620 96324 118621 96388
rect 118555 96323 118621 96324
rect 171363 80612 171429 80613
rect 171363 80548 171364 80612
rect 171428 80548 171429 80612
rect 171363 80547 171429 80548
rect 141003 80204 141069 80205
rect 141003 80140 141004 80204
rect 141068 80140 141069 80204
rect 141003 80139 141069 80140
rect 144867 80204 144933 80205
rect 144867 80140 144868 80204
rect 144932 80140 144933 80204
rect 144867 80139 144933 80140
rect 152411 80204 152477 80205
rect 152411 80140 152412 80204
rect 152476 80140 152477 80204
rect 152411 80139 152477 80140
rect 163451 80204 163517 80205
rect 163451 80140 163452 80204
rect 163516 80140 163517 80204
rect 163451 80139 163517 80140
rect 129779 80068 129845 80069
rect 129779 80004 129780 80068
rect 129844 80004 129845 80068
rect 129779 80003 129845 80004
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 126283 79932 126349 79933
rect 126283 79868 126284 79932
rect 126348 79868 126349 79932
rect 127387 79932 127453 79933
rect 127387 79930 127388 79932
rect 126283 79867 126349 79868
rect 127206 79870 127388 79930
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125915 77892 125981 77893
rect 125915 77828 125916 77892
rect 125980 77828 125981 77892
rect 125915 77827 125981 77828
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 125918 4861 125978 77827
rect 126286 77757 126346 79867
rect 126283 77756 126349 77757
rect 126283 77692 126284 77756
rect 126348 77692 126349 77756
rect 126283 77691 126349 77692
rect 127206 7581 127266 79870
rect 127387 79868 127388 79870
rect 127452 79868 127453 79932
rect 127755 79932 127821 79933
rect 127755 79930 127756 79932
rect 127387 79867 127453 79868
rect 127574 79870 127756 79930
rect 127387 79796 127453 79797
rect 127387 79732 127388 79796
rect 127452 79732 127453 79796
rect 127387 79731 127453 79732
rect 127203 7580 127269 7581
rect 127203 7516 127204 7580
rect 127268 7516 127269 7580
rect 127203 7515 127269 7516
rect 125915 4860 125981 4861
rect 125915 4796 125916 4860
rect 125980 4796 125981 4860
rect 125915 4795 125981 4796
rect 127390 3365 127450 79731
rect 127574 77893 127634 79870
rect 127755 79868 127756 79870
rect 127820 79868 127821 79932
rect 127755 79867 127821 79868
rect 128491 79932 128557 79933
rect 128491 79868 128492 79932
rect 128556 79868 128557 79932
rect 128491 79867 128557 79868
rect 129227 79932 129293 79933
rect 129227 79868 129228 79932
rect 129292 79868 129293 79932
rect 129227 79867 129293 79868
rect 127571 77892 127637 77893
rect 127571 77828 127572 77892
rect 127636 77828 127637 77892
rect 127571 77827 127637 77828
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127387 3364 127453 3365
rect 127387 3300 127388 3364
rect 127452 3300 127453 3364
rect 127387 3299 127453 3300
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 6930 128554 79867
rect 128675 79660 128741 79661
rect 128675 79596 128676 79660
rect 128740 79596 128741 79660
rect 128675 79595 128741 79596
rect 128678 8941 128738 79595
rect 128859 78844 128925 78845
rect 128859 78780 128860 78844
rect 128924 78780 128925 78844
rect 128859 78779 128925 78780
rect 128862 73813 128922 78779
rect 129230 78709 129290 79867
rect 129227 78708 129293 78709
rect 129227 78644 129228 78708
rect 129292 78644 129293 78708
rect 129227 78643 129293 78644
rect 128859 73812 128925 73813
rect 128859 73748 128860 73812
rect 128924 73748 128925 73812
rect 128859 73747 128925 73748
rect 129782 9077 129842 80003
rect 130883 79932 130949 79933
rect 130883 79868 130884 79932
rect 130948 79868 130949 79932
rect 130883 79867 130949 79868
rect 132171 79932 132237 79933
rect 132171 79868 132172 79932
rect 132236 79868 132237 79932
rect 132171 79867 132237 79868
rect 133459 79932 133525 79933
rect 133459 79868 133460 79932
rect 133524 79868 133525 79932
rect 133459 79867 133525 79868
rect 138059 79932 138125 79933
rect 138059 79868 138060 79932
rect 138124 79868 138125 79932
rect 138059 79867 138125 79868
rect 139163 79932 139229 79933
rect 139163 79868 139164 79932
rect 139228 79868 139229 79932
rect 139163 79867 139229 79868
rect 140635 79932 140701 79933
rect 140635 79868 140636 79932
rect 140700 79868 140701 79932
rect 140635 79867 140701 79868
rect 130331 79796 130397 79797
rect 130331 79732 130332 79796
rect 130396 79732 130397 79796
rect 130331 79731 130397 79732
rect 130147 78844 130213 78845
rect 130147 78780 130148 78844
rect 130212 78780 130213 78844
rect 130147 78779 130213 78780
rect 129963 78708 130029 78709
rect 129963 78644 129964 78708
rect 130028 78644 130029 78708
rect 129963 78643 130029 78644
rect 129966 9213 130026 78643
rect 130150 73949 130210 78779
rect 130334 74085 130394 79731
rect 130886 77310 130946 79867
rect 131251 79660 131317 79661
rect 131251 79596 131252 79660
rect 131316 79596 131317 79660
rect 131251 79595 131317 79596
rect 130886 77250 131130 77310
rect 131070 74221 131130 77250
rect 131067 74220 131133 74221
rect 131067 74156 131068 74220
rect 131132 74156 131133 74220
rect 131067 74155 131133 74156
rect 130331 74084 130397 74085
rect 130331 74020 130332 74084
rect 130396 74020 130397 74084
rect 130331 74019 130397 74020
rect 130147 73948 130213 73949
rect 130147 73884 130148 73948
rect 130212 73884 130213 73948
rect 130147 73883 130213 73884
rect 131254 10301 131314 79595
rect 131435 78708 131501 78709
rect 131435 78644 131436 78708
rect 131500 78644 131501 78708
rect 131435 78643 131501 78644
rect 131251 10300 131317 10301
rect 131251 10236 131252 10300
rect 131316 10236 131317 10300
rect 131251 10235 131317 10236
rect 129963 9212 130029 9213
rect 129963 9148 129964 9212
rect 130028 9148 130029 9212
rect 129963 9147 130029 9148
rect 129779 9076 129845 9077
rect 129779 9012 129780 9076
rect 129844 9012 129845 9076
rect 129779 9011 129845 9012
rect 128675 8940 128741 8941
rect 128675 8876 128676 8940
rect 128740 8876 128741 8940
rect 128675 8875 128741 8876
rect 128494 6870 128738 6930
rect 128678 6221 128738 6870
rect 131438 6357 131498 78643
rect 132174 78165 132234 79867
rect 133091 79660 133157 79661
rect 133091 79596 133092 79660
rect 133156 79596 133157 79660
rect 133091 79595 133157 79596
rect 132171 78164 132237 78165
rect 132171 78100 132172 78164
rect 132236 78100 132237 78164
rect 132171 78099 132237 78100
rect 131987 77756 132053 77757
rect 131987 77692 131988 77756
rect 132052 77692 132053 77756
rect 131987 77691 132053 77692
rect 131435 6356 131501 6357
rect 131435 6292 131436 6356
rect 131500 6292 131501 6356
rect 131435 6291 131501 6292
rect 128675 6220 128741 6221
rect 128675 6156 128676 6220
rect 128740 6156 128741 6220
rect 128675 6155 128741 6156
rect 131990 3773 132050 77691
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131987 3772 132053 3773
rect 131987 3708 131988 3772
rect 132052 3708 132053 3772
rect 131987 3707 132053 3708
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 10437 133154 79595
rect 133275 78028 133341 78029
rect 133275 77964 133276 78028
rect 133340 77964 133341 78028
rect 133275 77963 133341 77964
rect 133278 44845 133338 77963
rect 133462 77893 133522 79867
rect 135299 79796 135365 79797
rect 135299 79732 135300 79796
rect 135364 79732 135365 79796
rect 135299 79731 135365 79732
rect 137875 79796 137941 79797
rect 137875 79732 137876 79796
rect 137940 79732 137941 79796
rect 137875 79731 137941 79732
rect 134011 78708 134077 78709
rect 134011 78644 134012 78708
rect 134076 78644 134077 78708
rect 134011 78643 134077 78644
rect 133643 78300 133709 78301
rect 133643 78236 133644 78300
rect 133708 78236 133709 78300
rect 133643 78235 133709 78236
rect 133459 77892 133525 77893
rect 133459 77828 133460 77892
rect 133524 77828 133525 77892
rect 133459 77827 133525 77828
rect 133275 44844 133341 44845
rect 133275 44780 133276 44844
rect 133340 44780 133341 44844
rect 133275 44779 133341 44780
rect 133091 10436 133157 10437
rect 133091 10372 133092 10436
rect 133156 10372 133157 10436
rect 133091 10371 133157 10372
rect 133646 8805 133706 78235
rect 134014 10573 134074 78643
rect 134195 78028 134261 78029
rect 134195 77964 134196 78028
rect 134260 77964 134261 78028
rect 134195 77963 134261 77964
rect 134931 78028 134997 78029
rect 134931 77964 134932 78028
rect 134996 77964 134997 78028
rect 134931 77963 134997 77964
rect 134011 10572 134077 10573
rect 134011 10508 134012 10572
rect 134076 10508 134077 10572
rect 134011 10507 134077 10508
rect 133643 8804 133709 8805
rect 133643 8740 133644 8804
rect 133708 8740 133709 8804
rect 133643 8739 133709 8740
rect 134198 7717 134258 77963
rect 134934 17917 134994 77963
rect 135302 74493 135362 79731
rect 136403 78844 136469 78845
rect 136403 78780 136404 78844
rect 136468 78780 136469 78844
rect 136403 78779 136469 78780
rect 137691 78844 137757 78845
rect 137691 78780 137692 78844
rect 137756 78780 137757 78844
rect 137691 78779 137757 78780
rect 136035 77892 136101 77893
rect 136035 77828 136036 77892
rect 136100 77828 136101 77892
rect 136035 77827 136101 77828
rect 135299 74492 135365 74493
rect 135299 74428 135300 74492
rect 135364 74428 135365 74492
rect 135299 74427 135365 74428
rect 134931 17916 134997 17917
rect 134931 17852 134932 17916
rect 134996 17852 134997 17916
rect 134931 17851 134997 17852
rect 136038 17645 136098 77827
rect 136219 77076 136285 77077
rect 136219 77012 136220 77076
rect 136284 77012 136285 77076
rect 136219 77011 136285 77012
rect 136035 17644 136101 17645
rect 136035 17580 136036 17644
rect 136100 17580 136101 17644
rect 136035 17579 136101 17580
rect 134195 7716 134261 7717
rect 134195 7652 134196 7716
rect 134260 7652 134261 7716
rect 134195 7651 134261 7652
rect 136222 3637 136282 77011
rect 136406 4045 136466 78779
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 4044 136469 4045
rect 136403 3980 136404 4044
rect 136468 3980 136469 4044
rect 136403 3979 136469 3980
rect 136219 3636 136285 3637
rect 136219 3572 136220 3636
rect 136284 3572 136285 3636
rect 136219 3571 136285 3572
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137694 6221 137754 78779
rect 137691 6220 137757 6221
rect 137691 6156 137692 6220
rect 137756 6156 137757 6220
rect 137691 6155 137757 6156
rect 137878 4861 137938 79731
rect 138062 78709 138122 79867
rect 138979 79796 139045 79797
rect 138979 79732 138980 79796
rect 139044 79732 139045 79796
rect 138979 79731 139045 79732
rect 138611 79660 138677 79661
rect 138611 79596 138612 79660
rect 138676 79596 138677 79660
rect 138611 79595 138677 79596
rect 138059 78708 138125 78709
rect 138059 78644 138060 78708
rect 138124 78644 138125 78708
rect 138059 78643 138125 78644
rect 138059 77892 138125 77893
rect 138059 77828 138060 77892
rect 138124 77828 138125 77892
rect 138059 77827 138125 77828
rect 138062 77349 138122 77827
rect 138059 77348 138125 77349
rect 138059 77284 138060 77348
rect 138124 77284 138125 77348
rect 138059 77283 138125 77284
rect 138614 61437 138674 79595
rect 138795 78708 138861 78709
rect 138795 78644 138796 78708
rect 138860 78644 138861 78708
rect 138795 78643 138861 78644
rect 138798 69597 138858 78643
rect 138795 69596 138861 69597
rect 138795 69532 138796 69596
rect 138860 69532 138861 69596
rect 138795 69531 138861 69532
rect 138982 62797 139042 79731
rect 139166 75717 139226 79867
rect 139531 79660 139597 79661
rect 139531 79596 139532 79660
rect 139596 79596 139597 79660
rect 139531 79595 139597 79596
rect 139534 75989 139594 79595
rect 140451 78844 140517 78845
rect 140451 78780 140452 78844
rect 140516 78780 140517 78844
rect 140451 78779 140517 78780
rect 139531 75988 139597 75989
rect 139531 75924 139532 75988
rect 139596 75924 139597 75988
rect 139531 75923 139597 75924
rect 140083 75852 140149 75853
rect 140083 75788 140084 75852
rect 140148 75788 140149 75852
rect 140083 75787 140149 75788
rect 139163 75716 139229 75717
rect 139163 75652 139164 75716
rect 139228 75652 139229 75716
rect 139163 75651 139229 75652
rect 138979 62796 139045 62797
rect 138979 62732 138980 62796
rect 139044 62732 139045 62796
rect 138979 62731 139045 62732
rect 138611 61436 138677 61437
rect 138611 61372 138612 61436
rect 138676 61372 138677 61436
rect 138611 61371 138677 61372
rect 140086 6085 140146 75787
rect 140267 73132 140333 73133
rect 140267 73068 140268 73132
rect 140332 73068 140333 73132
rect 140267 73067 140333 73068
rect 140270 65517 140330 73067
rect 140267 65516 140333 65517
rect 140267 65452 140268 65516
rect 140332 65452 140333 65516
rect 140267 65451 140333 65452
rect 140454 17101 140514 78779
rect 140638 78301 140698 79867
rect 140635 78300 140701 78301
rect 140635 78236 140636 78300
rect 140700 78236 140701 78300
rect 140635 78235 140701 78236
rect 141006 34101 141066 80139
rect 143211 79932 143277 79933
rect 143211 79868 143212 79932
rect 143276 79868 143277 79932
rect 143211 79867 143277 79868
rect 144131 79932 144197 79933
rect 144131 79868 144132 79932
rect 144196 79868 144197 79932
rect 144131 79867 144197 79868
rect 144683 79932 144749 79933
rect 144683 79868 144684 79932
rect 144748 79868 144749 79932
rect 144683 79867 144749 79868
rect 141371 79796 141437 79797
rect 141371 79732 141372 79796
rect 141436 79732 141437 79796
rect 141371 79731 141437 79732
rect 142843 79796 142909 79797
rect 142843 79732 142844 79796
rect 142908 79732 142909 79796
rect 142843 79731 142909 79732
rect 141374 78165 141434 79731
rect 141371 78164 141437 78165
rect 141371 78100 141372 78164
rect 141436 78100 141437 78164
rect 141371 78099 141437 78100
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 34100 141069 34101
rect 141003 34036 141004 34100
rect 141068 34036 141069 34100
rect 141003 34035 141069 34036
rect 140451 17100 140517 17101
rect 140451 17036 140452 17100
rect 140516 17036 140517 17100
rect 140451 17035 140517 17036
rect 140083 6084 140149 6085
rect 140083 6020 140084 6084
rect 140148 6020 140149 6084
rect 140083 6019 140149 6020
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 6901 142906 79731
rect 143027 76668 143093 76669
rect 143027 76604 143028 76668
rect 143092 76604 143093 76668
rect 143027 76603 143093 76604
rect 143030 33965 143090 76603
rect 143027 33964 143093 33965
rect 143027 33900 143028 33964
rect 143092 33900 143093 33964
rect 143027 33899 143093 33900
rect 143214 13293 143274 79867
rect 144134 76669 144194 79867
rect 144315 79796 144381 79797
rect 144315 79732 144316 79796
rect 144380 79732 144381 79796
rect 144315 79731 144381 79732
rect 144499 79796 144565 79797
rect 144499 79732 144500 79796
rect 144564 79732 144565 79796
rect 144499 79731 144565 79732
rect 144131 76668 144197 76669
rect 144131 76604 144132 76668
rect 144196 76604 144197 76668
rect 144131 76603 144197 76604
rect 144318 27029 144378 79731
rect 144315 27028 144381 27029
rect 144315 26964 144316 27028
rect 144380 26964 144381 27028
rect 144315 26963 144381 26964
rect 144502 20501 144562 79731
rect 144499 20500 144565 20501
rect 144499 20436 144500 20500
rect 144564 20436 144565 20500
rect 144499 20435 144565 20436
rect 143211 13292 143277 13293
rect 143211 13228 143212 13292
rect 143276 13228 143277 13292
rect 143211 13227 143277 13228
rect 142843 6900 142909 6901
rect 142843 6836 142844 6900
rect 142908 6836 142909 6900
rect 142843 6835 142909 6836
rect 144686 6765 144746 79867
rect 144870 76261 144930 80139
rect 145419 80068 145485 80069
rect 145419 80004 145420 80068
rect 145484 80004 145485 80068
rect 145419 80003 145485 80004
rect 145051 79932 145117 79933
rect 145051 79868 145052 79932
rect 145116 79868 145117 79932
rect 145051 79867 145117 79868
rect 144867 76260 144933 76261
rect 144867 76196 144868 76260
rect 144932 76196 144933 76260
rect 144867 76195 144933 76196
rect 145054 75989 145114 79867
rect 145422 79661 145482 80003
rect 147075 79932 147141 79933
rect 147075 79868 147076 79932
rect 147140 79868 147141 79932
rect 147075 79867 147141 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148179 79867 148245 79868
rect 148731 79932 148797 79933
rect 148731 79868 148732 79932
rect 148796 79868 148797 79932
rect 148731 79867 148797 79868
rect 149651 79932 149717 79933
rect 149651 79868 149652 79932
rect 149716 79868 149717 79932
rect 149651 79867 149717 79868
rect 150571 79932 150637 79933
rect 150571 79868 150572 79932
rect 150636 79868 150637 79932
rect 150571 79867 150637 79868
rect 151859 79932 151925 79933
rect 151859 79868 151860 79932
rect 151924 79868 151925 79932
rect 151859 79867 151925 79868
rect 145603 79796 145669 79797
rect 145603 79732 145604 79796
rect 145668 79732 145669 79796
rect 145603 79731 145669 79732
rect 145419 79660 145485 79661
rect 145419 79596 145420 79660
rect 145484 79596 145485 79660
rect 145419 79595 145485 79596
rect 145051 75988 145117 75989
rect 145051 75924 145052 75988
rect 145116 75924 145117 75988
rect 145051 75923 145117 75924
rect 145419 75852 145485 75853
rect 145419 75788 145420 75852
rect 145484 75788 145485 75852
rect 145419 75787 145485 75788
rect 145235 74220 145301 74221
rect 145235 74156 145236 74220
rect 145300 74156 145301 74220
rect 145235 74155 145301 74156
rect 145238 33829 145298 74155
rect 145235 33828 145301 33829
rect 145235 33764 145236 33828
rect 145300 33764 145301 33828
rect 145235 33763 145301 33764
rect 145422 14925 145482 75787
rect 145419 14924 145485 14925
rect 145419 14860 145420 14924
rect 145484 14860 145485 14924
rect 145419 14859 145485 14860
rect 144683 6764 144749 6765
rect 144683 6700 144684 6764
rect 144748 6700 144749 6764
rect 144683 6699 144749 6700
rect 145606 6629 145666 79731
rect 145794 75454 146414 78000
rect 146891 75988 146957 75989
rect 146891 75924 146892 75988
rect 146956 75924 146957 75988
rect 146891 75923 146957 75924
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 6628 145669 6629
rect 145603 6564 145604 6628
rect 145668 6564 145669 6628
rect 145603 6563 145669 6564
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 146894 9621 146954 75923
rect 147078 17781 147138 79867
rect 147259 79796 147325 79797
rect 147259 79732 147260 79796
rect 147324 79732 147325 79796
rect 147259 79731 147325 79732
rect 147075 17780 147141 17781
rect 147075 17716 147076 17780
rect 147140 17716 147141 17780
rect 147075 17715 147141 17716
rect 147262 14789 147322 79731
rect 148182 76669 148242 79867
rect 148547 79796 148613 79797
rect 148547 79732 148548 79796
rect 148612 79732 148613 79796
rect 148547 79731 148613 79732
rect 148363 76804 148429 76805
rect 148363 76740 148364 76804
rect 148428 76740 148429 76804
rect 148363 76739 148429 76740
rect 148179 76668 148245 76669
rect 148179 76604 148180 76668
rect 148244 76604 148245 76668
rect 148179 76603 148245 76604
rect 147259 14788 147325 14789
rect 147259 14724 147260 14788
rect 147324 14724 147325 14788
rect 147259 14723 147325 14724
rect 146891 9620 146957 9621
rect 146891 9556 146892 9620
rect 146956 9556 146957 9620
rect 146891 9555 146957 9556
rect 148366 6493 148426 76739
rect 148550 17509 148610 79731
rect 148547 17508 148613 17509
rect 148547 17444 148548 17508
rect 148612 17444 148613 17508
rect 148547 17443 148613 17444
rect 148734 9485 148794 79867
rect 149467 77348 149533 77349
rect 149467 77284 149468 77348
rect 149532 77284 149533 77348
rect 149467 77283 149533 77284
rect 148915 76668 148981 76669
rect 148915 76604 148916 76668
rect 148980 76604 148981 76668
rect 148915 76603 148981 76604
rect 148918 72589 148978 76603
rect 148915 72588 148981 72589
rect 148915 72524 148916 72588
rect 148980 72524 148981 72588
rect 148915 72523 148981 72524
rect 149470 35325 149530 77283
rect 149467 35324 149533 35325
rect 149467 35260 149468 35324
rect 149532 35260 149533 35324
rect 149467 35259 149533 35260
rect 149654 26893 149714 79867
rect 150019 79796 150085 79797
rect 150019 79732 150020 79796
rect 150084 79732 150085 79796
rect 150019 79731 150085 79732
rect 149835 78164 149901 78165
rect 149835 78100 149836 78164
rect 149900 78100 149901 78164
rect 149835 78099 149901 78100
rect 149651 26892 149717 26893
rect 149651 26828 149652 26892
rect 149716 26828 149717 26892
rect 149651 26827 149717 26828
rect 148731 9484 148797 9485
rect 148731 9420 148732 9484
rect 148796 9420 148797 9484
rect 148731 9419 148797 9420
rect 149838 9349 149898 78099
rect 149835 9348 149901 9349
rect 149835 9284 149836 9348
rect 149900 9284 149901 9348
rect 149835 9283 149901 9284
rect 150022 9213 150082 79731
rect 150574 78165 150634 79867
rect 151491 79660 151557 79661
rect 151491 79596 151492 79660
rect 151556 79596 151557 79660
rect 151491 79595 151557 79596
rect 151307 78844 151373 78845
rect 151307 78780 151308 78844
rect 151372 78780 151373 78844
rect 151307 78779 151373 78780
rect 150571 78164 150637 78165
rect 150571 78100 150572 78164
rect 150636 78100 150637 78164
rect 150571 78099 150637 78100
rect 150294 43954 150914 78000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150019 9212 150085 9213
rect 150019 9148 150020 9212
rect 150084 9148 150085 9212
rect 150019 9147 150085 9148
rect 150294 7954 150914 43398
rect 151310 31109 151370 78779
rect 151307 31108 151373 31109
rect 151307 31044 151308 31108
rect 151372 31044 151373 31108
rect 151307 31043 151373 31044
rect 151494 28389 151554 79595
rect 151862 78709 151922 79867
rect 151675 78708 151741 78709
rect 151675 78644 151676 78708
rect 151740 78644 151741 78708
rect 151675 78643 151741 78644
rect 151859 78708 151925 78709
rect 151859 78644 151860 78708
rect 151924 78644 151925 78708
rect 151859 78643 151925 78644
rect 151491 28388 151557 28389
rect 151491 28324 151492 28388
rect 151556 28324 151557 28388
rect 151491 28323 151557 28324
rect 151678 12069 151738 78643
rect 151675 12068 151741 12069
rect 151675 12004 151676 12068
rect 151740 12004 151741 12068
rect 151675 12003 151741 12004
rect 152414 9077 152474 80139
rect 153147 79932 153213 79933
rect 153147 79868 153148 79932
rect 153212 79868 153213 79932
rect 153147 79867 153213 79868
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 153883 79867 153949 79868
rect 155723 79932 155789 79933
rect 155723 79868 155724 79932
rect 155788 79868 155789 79932
rect 155723 79867 155789 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79930 156893 79932
rect 157931 79932 157997 79933
rect 156892 79870 157074 79930
rect 156892 79868 156893 79870
rect 156827 79867 156893 79868
rect 152779 79796 152845 79797
rect 152779 79732 152780 79796
rect 152844 79732 152845 79796
rect 152779 79731 152845 79732
rect 152595 77348 152661 77349
rect 152595 77284 152596 77348
rect 152660 77284 152661 77348
rect 152595 77283 152661 77284
rect 152598 68237 152658 77283
rect 152595 68236 152661 68237
rect 152595 68172 152596 68236
rect 152660 68172 152661 68236
rect 152595 68171 152661 68172
rect 152782 51781 152842 79731
rect 153150 77077 153210 79867
rect 153147 77076 153213 77077
rect 153147 77012 153148 77076
rect 153212 77012 153213 77076
rect 153147 77011 153213 77012
rect 153886 58581 153946 79867
rect 154067 79796 154133 79797
rect 154067 79732 154068 79796
rect 154132 79732 154133 79796
rect 154067 79731 154133 79732
rect 154435 79796 154501 79797
rect 154435 79732 154436 79796
rect 154500 79732 154501 79796
rect 154435 79731 154501 79732
rect 153883 58580 153949 58581
rect 153883 58516 153884 58580
rect 153948 58516 153949 58580
rect 153883 58515 153949 58516
rect 152779 51780 152845 51781
rect 152779 51716 152780 51780
rect 152844 51716 152845 51780
rect 152779 51715 152845 51716
rect 154070 16149 154130 79731
rect 154251 79660 154317 79661
rect 154251 79596 154252 79660
rect 154316 79596 154317 79660
rect 154251 79595 154317 79596
rect 154067 16148 154133 16149
rect 154067 16084 154068 16148
rect 154132 16084 154133 16148
rect 154067 16083 154133 16084
rect 154254 14653 154314 79595
rect 154251 14652 154317 14653
rect 154251 14588 154252 14652
rect 154316 14588 154317 14652
rect 154251 14587 154317 14588
rect 154438 13157 154498 79731
rect 154794 48454 155414 78000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13156 154501 13157
rect 154435 13092 154436 13156
rect 154500 13092 154501 13156
rect 154435 13091 154501 13092
rect 154794 12454 155414 47898
rect 155726 16013 155786 79867
rect 156827 79660 156893 79661
rect 156827 79596 156828 79660
rect 156892 79596 156893 79660
rect 156827 79595 156893 79596
rect 156643 78708 156709 78709
rect 156643 78644 156644 78708
rect 156708 78644 156709 78708
rect 156643 78643 156709 78644
rect 155723 16012 155789 16013
rect 155723 15948 155724 16012
rect 155788 15948 155789 16012
rect 155723 15947 155789 15948
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 152411 9076 152477 9077
rect 152411 9012 152412 9076
rect 152476 9012 152477 9076
rect 152411 9011 152477 9012
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 148363 6492 148429 6493
rect 148363 6428 148364 6492
rect 148428 6428 148429 6492
rect 148363 6427 148429 6428
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 156646 8941 156706 78643
rect 156830 20365 156890 79595
rect 156827 20364 156893 20365
rect 156827 20300 156828 20364
rect 156892 20300 156893 20364
rect 156827 20299 156893 20300
rect 157014 17373 157074 79870
rect 157931 79868 157932 79932
rect 157996 79868 157997 79932
rect 157931 79867 157997 79868
rect 158299 79932 158365 79933
rect 158299 79868 158300 79932
rect 158364 79930 158365 79932
rect 159955 79932 160021 79933
rect 158364 79870 158546 79930
rect 158364 79868 158365 79870
rect 158299 79867 158365 79868
rect 157747 79660 157813 79661
rect 157747 79596 157748 79660
rect 157812 79596 157813 79660
rect 157747 79595 157813 79596
rect 157750 77349 157810 79595
rect 157934 77893 157994 79867
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 157931 77892 157997 77893
rect 157931 77828 157932 77892
rect 157996 77828 157997 77892
rect 157931 77827 157997 77828
rect 157747 77348 157813 77349
rect 157747 77284 157748 77348
rect 157812 77284 157813 77348
rect 157747 77283 157813 77284
rect 157931 76668 157997 76669
rect 157931 76604 157932 76668
rect 157996 76604 157997 76668
rect 157931 76603 157997 76604
rect 157934 29613 157994 76603
rect 158115 74492 158181 74493
rect 158115 74428 158116 74492
rect 158180 74428 158181 74492
rect 158115 74427 158181 74428
rect 157931 29612 157997 29613
rect 157931 29548 157932 29612
rect 157996 29548 157997 29612
rect 157931 29547 157997 29548
rect 157011 17372 157077 17373
rect 157011 17308 157012 17372
rect 157076 17308 157077 17372
rect 157011 17307 157077 17308
rect 158118 17237 158178 74427
rect 158115 17236 158181 17237
rect 158115 17172 158116 17236
rect 158180 17172 158181 17236
rect 158115 17171 158181 17172
rect 158302 11933 158362 79731
rect 158299 11932 158365 11933
rect 158299 11868 158300 11932
rect 158364 11868 158365 11932
rect 158299 11867 158365 11868
rect 158486 10301 158546 79870
rect 159955 79868 159956 79932
rect 160020 79868 160021 79932
rect 159955 79867 160021 79868
rect 160875 79932 160941 79933
rect 160875 79868 160876 79932
rect 160940 79868 160941 79932
rect 160875 79867 160941 79868
rect 161059 79932 161125 79933
rect 161059 79868 161060 79932
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 161427 79932 161493 79933
rect 161427 79868 161428 79932
rect 161492 79868 161493 79932
rect 161427 79867 161493 79868
rect 161795 79932 161861 79933
rect 161795 79868 161796 79932
rect 161860 79868 161861 79932
rect 161795 79867 161861 79868
rect 159958 78845 160018 79867
rect 160507 79796 160573 79797
rect 160507 79732 160508 79796
rect 160572 79732 160573 79796
rect 160507 79731 160573 79732
rect 160323 79660 160389 79661
rect 160323 79596 160324 79660
rect 160388 79596 160389 79660
rect 160323 79595 160389 79596
rect 159955 78844 160021 78845
rect 159955 78780 159956 78844
rect 160020 78780 160021 78844
rect 159955 78779 160021 78780
rect 160326 78709 160386 79595
rect 160323 78708 160389 78709
rect 160323 78644 160324 78708
rect 160388 78644 160389 78708
rect 160323 78643 160389 78644
rect 159035 75988 159101 75989
rect 159035 75924 159036 75988
rect 159100 75924 159101 75988
rect 159035 75923 159101 75924
rect 159038 21317 159098 75923
rect 159294 52954 159914 78000
rect 160510 75989 160570 79731
rect 160691 79660 160757 79661
rect 160691 79596 160692 79660
rect 160756 79596 160757 79660
rect 160691 79595 160757 79596
rect 160507 75988 160573 75989
rect 160507 75924 160508 75988
rect 160572 75924 160573 75988
rect 160507 75923 160573 75924
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 21316 159101 21317
rect 159035 21252 159036 21316
rect 159100 21252 159101 21316
rect 159035 21251 159101 21252
rect 159294 16954 159914 52398
rect 160694 20093 160754 79595
rect 160878 75853 160938 79867
rect 160875 75852 160941 75853
rect 160875 75788 160876 75852
rect 160940 75788 160941 75852
rect 160875 75787 160941 75788
rect 161062 20229 161122 79867
rect 161430 75037 161490 79867
rect 161798 75853 161858 79867
rect 162715 79796 162781 79797
rect 162715 79732 162716 79796
rect 162780 79732 162781 79796
rect 162715 79731 162781 79732
rect 163083 79796 163149 79797
rect 163083 79732 163084 79796
rect 163148 79732 163149 79796
rect 163083 79731 163149 79732
rect 162531 79660 162597 79661
rect 162531 79596 162532 79660
rect 162596 79596 162597 79660
rect 162531 79595 162597 79596
rect 162347 75988 162413 75989
rect 162347 75924 162348 75988
rect 162412 75924 162413 75988
rect 162347 75923 162413 75924
rect 161795 75852 161861 75853
rect 161795 75788 161796 75852
rect 161860 75788 161861 75852
rect 161795 75787 161861 75788
rect 161427 75036 161493 75037
rect 161427 74972 161428 75036
rect 161492 74972 161493 75036
rect 161427 74971 161493 74972
rect 162350 22813 162410 75923
rect 162347 22812 162413 22813
rect 162347 22748 162348 22812
rect 162412 22748 162413 22812
rect 162347 22747 162413 22748
rect 161059 20228 161125 20229
rect 161059 20164 161060 20228
rect 161124 20164 161125 20228
rect 161059 20163 161125 20164
rect 160691 20092 160757 20093
rect 160691 20028 160692 20092
rect 160756 20028 160757 20092
rect 160691 20027 160757 20028
rect 162534 19957 162594 79595
rect 162531 19956 162597 19957
rect 162531 19892 162532 19956
rect 162596 19892 162597 19956
rect 162531 19891 162597 19892
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 10300 158549 10301
rect 158483 10236 158484 10300
rect 158548 10236 158549 10300
rect 158483 10235 158549 10236
rect 156643 8940 156709 8941
rect 156643 8876 156644 8940
rect 156708 8876 156709 8940
rect 156643 8875 156709 8876
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 162718 15877 162778 79731
rect 163086 77349 163146 79731
rect 163267 79660 163333 79661
rect 163267 79596 163268 79660
rect 163332 79596 163333 79660
rect 163267 79595 163333 79596
rect 163270 78709 163330 79595
rect 163267 78708 163333 78709
rect 163267 78644 163268 78708
rect 163332 78644 163333 78708
rect 163267 78643 163333 78644
rect 163083 77348 163149 77349
rect 163083 77284 163084 77348
rect 163148 77284 163149 77348
rect 163083 77283 163149 77284
rect 163454 35189 163514 80139
rect 171366 79933 171426 80547
rect 172283 80340 172349 80341
rect 172283 80276 172284 80340
rect 172348 80276 172349 80340
rect 172283 80275 172349 80276
rect 172099 80204 172165 80205
rect 172099 80140 172100 80204
rect 172164 80140 172165 80204
rect 172099 80139 172165 80140
rect 165475 79932 165541 79933
rect 165475 79868 165476 79932
rect 165540 79868 165541 79932
rect 165475 79867 165541 79868
rect 166027 79932 166093 79933
rect 166027 79868 166028 79932
rect 166092 79868 166093 79932
rect 166027 79867 166093 79868
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 167315 79932 167381 79933
rect 167315 79868 167316 79932
rect 167380 79868 167381 79932
rect 168051 79932 168117 79933
rect 168051 79930 168052 79932
rect 167315 79867 167381 79868
rect 167870 79870 168052 79930
rect 163635 79660 163701 79661
rect 163635 79596 163636 79660
rect 163700 79596 163701 79660
rect 163635 79595 163701 79596
rect 163451 35188 163517 35189
rect 163451 35124 163452 35188
rect 163516 35124 163517 35188
rect 163451 35123 163517 35124
rect 162715 15876 162781 15877
rect 162715 15812 162716 15876
rect 162780 15812 162781 15876
rect 162715 15811 162781 15812
rect 163638 5133 163698 79595
rect 165107 78844 165173 78845
rect 165107 78780 165108 78844
rect 165172 78780 165173 78844
rect 165107 78779 165173 78780
rect 163794 57454 164414 78000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 165110 55861 165170 78779
rect 165291 75988 165357 75989
rect 165291 75924 165292 75988
rect 165356 75924 165357 75988
rect 165291 75923 165357 75924
rect 165107 55860 165173 55861
rect 165107 55796 165108 55860
rect 165172 55796 165173 55860
rect 165107 55795 165173 55796
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 5132 163701 5133
rect 163635 5068 163636 5132
rect 163700 5068 163701 5132
rect 163635 5067 163701 5068
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 165294 14517 165354 75923
rect 165291 14516 165357 14517
rect 165291 14452 165292 14516
rect 165356 14452 165357 14516
rect 165291 14451 165357 14452
rect 165478 11797 165538 79867
rect 166030 75989 166090 79867
rect 166214 75989 166274 79867
rect 166395 79796 166461 79797
rect 166395 79732 166396 79796
rect 166460 79732 166461 79796
rect 166395 79731 166461 79732
rect 166027 75988 166093 75989
rect 166027 75924 166028 75988
rect 166092 75924 166093 75988
rect 166027 75923 166093 75924
rect 166211 75988 166277 75989
rect 166211 75924 166212 75988
rect 166276 75924 166277 75988
rect 166211 75923 166277 75924
rect 166211 73268 166277 73269
rect 166211 73204 166212 73268
rect 166276 73204 166277 73268
rect 166211 73203 166277 73204
rect 166214 66877 166274 73203
rect 166211 66876 166277 66877
rect 166211 66812 166212 66876
rect 166276 66812 166277 66876
rect 166211 66811 166277 66812
rect 166398 28253 166458 79731
rect 166579 79660 166645 79661
rect 166579 79596 166580 79660
rect 166644 79596 166645 79660
rect 166579 79595 166645 79596
rect 166395 28252 166461 28253
rect 166395 28188 166396 28252
rect 166460 28188 166461 28252
rect 166395 28187 166461 28188
rect 166582 18733 166642 79595
rect 166763 76124 166829 76125
rect 166763 76060 166764 76124
rect 166828 76060 166829 76124
rect 166763 76059 166829 76060
rect 166579 18732 166645 18733
rect 166579 18668 166580 18732
rect 166644 18668 166645 18732
rect 166579 18667 166645 18668
rect 166766 13021 166826 76059
rect 167318 75989 167378 79867
rect 167683 79796 167749 79797
rect 167683 79732 167684 79796
rect 167748 79732 167749 79796
rect 167683 79731 167749 79732
rect 167315 75988 167381 75989
rect 167315 75924 167316 75988
rect 167380 75924 167381 75988
rect 167315 75923 167381 75924
rect 167686 18597 167746 79731
rect 167683 18596 167749 18597
rect 167683 18532 167684 18596
rect 167748 18532 167749 18596
rect 167683 18531 167749 18532
rect 166763 13020 166829 13021
rect 166763 12956 166764 13020
rect 166828 12956 166829 13020
rect 166763 12955 166829 12956
rect 165475 11796 165541 11797
rect 165475 11732 165476 11796
rect 165540 11732 165541 11796
rect 165475 11731 165541 11732
rect 167870 6357 167930 79870
rect 168051 79868 168052 79870
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 169891 79932 169957 79933
rect 169891 79868 169892 79932
rect 169956 79868 169957 79932
rect 169891 79867 169957 79868
rect 170811 79932 170877 79933
rect 170811 79868 170812 79932
rect 170876 79930 170877 79932
rect 171363 79932 171429 79933
rect 170876 79870 171058 79930
rect 170876 79868 170877 79870
rect 170811 79867 170877 79868
rect 169523 79660 169589 79661
rect 169523 79596 169524 79660
rect 169588 79596 169589 79660
rect 169523 79595 169589 79596
rect 168051 77484 168117 77485
rect 168051 77420 168052 77484
rect 168116 77420 168117 77484
rect 168051 77419 168117 77420
rect 167867 6356 167933 6357
rect 167867 6292 167868 6356
rect 167932 6292 167933 6356
rect 167867 6291 167933 6292
rect 168054 4997 168114 77419
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169526 30973 169586 79595
rect 169894 77485 169954 79867
rect 170627 79796 170693 79797
rect 170627 79732 170628 79796
rect 170692 79732 170693 79796
rect 170627 79731 170693 79732
rect 169891 77484 169957 77485
rect 169891 77420 169892 77484
rect 169956 77420 169957 77484
rect 169891 77419 169957 77420
rect 170443 77484 170509 77485
rect 170443 77420 170444 77484
rect 170508 77420 170509 77484
rect 170443 77419 170509 77420
rect 170446 73813 170506 77419
rect 170443 73812 170509 73813
rect 170443 73748 170444 73812
rect 170508 73748 170509 73812
rect 170443 73747 170509 73748
rect 169523 30972 169589 30973
rect 169523 30908 169524 30972
rect 169588 30908 169589 30972
rect 169523 30907 169589 30908
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 4996 168117 4997
rect 168051 4932 168052 4996
rect 168116 4932 168117 4996
rect 168051 4931 168117 4932
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170630 22677 170690 79731
rect 170811 77348 170877 77349
rect 170811 77284 170812 77348
rect 170876 77284 170877 77348
rect 170811 77283 170877 77284
rect 170627 22676 170693 22677
rect 170627 22612 170628 22676
rect 170692 22612 170693 22676
rect 170627 22611 170693 22612
rect 170814 6221 170874 77283
rect 170811 6220 170877 6221
rect 170811 6156 170812 6220
rect 170876 6156 170877 6220
rect 170811 6155 170877 6156
rect 170998 4861 171058 79870
rect 171363 79868 171364 79932
rect 171428 79868 171429 79932
rect 171363 79867 171429 79868
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 171915 79867 171981 79868
rect 171918 79525 171978 79867
rect 171915 79524 171981 79525
rect 171915 79460 171916 79524
rect 171980 79460 171981 79524
rect 171915 79459 171981 79460
rect 171731 76260 171797 76261
rect 171731 76196 171732 76260
rect 171796 76196 171797 76260
rect 171731 76195 171797 76196
rect 170995 4860 171061 4861
rect 170995 4796 170996 4860
rect 171060 4796 171061 4860
rect 170995 4795 171061 4796
rect 171734 3365 171794 76195
rect 171915 75036 171981 75037
rect 171915 74972 171916 75036
rect 171980 74972 171981 75036
rect 171915 74971 171981 74972
rect 171918 3501 171978 74971
rect 172102 42125 172162 80139
rect 172286 72453 172346 80275
rect 173019 80204 173085 80205
rect 173019 80140 173020 80204
rect 173084 80202 173085 80204
rect 173084 80142 173266 80202
rect 173084 80140 173085 80142
rect 173019 80139 173085 80140
rect 172651 79932 172717 79933
rect 172651 79868 172652 79932
rect 172716 79930 172717 79932
rect 173019 79932 173085 79933
rect 172716 79870 172898 79930
rect 172716 79868 172717 79870
rect 172651 79867 172717 79868
rect 172651 79796 172717 79797
rect 172651 79732 172652 79796
rect 172716 79732 172717 79796
rect 172651 79731 172717 79732
rect 172654 79525 172714 79731
rect 172651 79524 172717 79525
rect 172651 79460 172652 79524
rect 172716 79460 172717 79524
rect 172651 79459 172717 79460
rect 172838 78845 172898 79870
rect 173019 79868 173020 79932
rect 173084 79868 173085 79932
rect 173019 79867 173085 79868
rect 172835 78844 172901 78845
rect 172835 78780 172836 78844
rect 172900 78780 172901 78844
rect 172835 78779 172901 78780
rect 173022 78709 173082 79867
rect 173206 78709 173266 80142
rect 186294 79954 186914 115398
rect 173387 79932 173453 79933
rect 173387 79868 173388 79932
rect 173452 79868 173453 79932
rect 173387 79867 173453 79868
rect 173939 79932 174005 79933
rect 173939 79868 173940 79932
rect 174004 79868 174005 79932
rect 173939 79867 174005 79868
rect 173390 79253 173450 79867
rect 173571 79796 173637 79797
rect 173571 79732 173572 79796
rect 173636 79732 173637 79796
rect 173571 79731 173637 79732
rect 173387 79252 173453 79253
rect 173387 79188 173388 79252
rect 173452 79188 173453 79252
rect 173387 79187 173453 79188
rect 173019 78708 173085 78709
rect 173019 78644 173020 78708
rect 173084 78644 173085 78708
rect 173019 78643 173085 78644
rect 173203 78708 173269 78709
rect 173203 78644 173204 78708
rect 173268 78644 173269 78708
rect 173203 78643 173269 78644
rect 173574 78573 173634 79731
rect 173571 78572 173637 78573
rect 173571 78508 173572 78572
rect 173636 78508 173637 78572
rect 173571 78507 173637 78508
rect 173942 78437 174002 79867
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 173939 78436 174005 78437
rect 173939 78372 173940 78436
rect 174004 78372 174005 78436
rect 173939 78371 174005 78372
rect 172283 72452 172349 72453
rect 172283 72388 172284 72452
rect 172348 72388 172349 72452
rect 172283 72387 172349 72388
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172099 42124 172165 42125
rect 172099 42060 172100 42124
rect 172164 42060 172165 42124
rect 172099 42059 172165 42060
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 171915 3500 171981 3501
rect 171915 3436 171916 3500
rect 171980 3436 171981 3500
rect 171915 3435 171981 3436
rect 171731 3364 171797 3365
rect 171731 3300 171732 3364
rect 171796 3300 171797 3364
rect 171731 3299 171797 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 172794 142000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew ground bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
